
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity controller_rom2 is
generic
	(
		ADDR_WIDTH : integer := 15 -- Specify your actual ROM size to save LEs and unnecessary block RAM usage.
	);
port (
	clk : in std_logic;
	reset_n : in std_logic := '1';
	addr : in std_logic_vector(ADDR_WIDTH-1 downto 0);
	q : out std_logic_vector(31 downto 0);
	-- Allow writes - defaults supplied to simplify projects that don't need to write.
	d : in std_logic_vector(31 downto 0) := X"00000000";
	we : in std_logic := '0';
	bytesel : in std_logic_vector(3 downto 0) := "1111"
);
end entity;

architecture rtl of controller_rom2 is

	signal addr1 : integer range 0 to 2**ADDR_WIDTH-1;

	--  build up 2D array to hold the memory
	type word_t is array (0 to 3) of std_logic_vector(7 downto 0);
	type ram_t is array (0 to 2 ** ADDR_WIDTH - 1) of word_t;

	signal ram : ram_t:=
	(

     0 => (x"4c",x"55",x"41",x"46"),
     1 => (x"00",x"30",x"3d",x"54"),
     2 => (x"00",x"00",x"1f",x"ef"),
     3 => (x"00",x"00",x"1f",x"f5"),
     4 => (x"00",x"00",x"1f",x"f9"),
     5 => (x"00",x"00",x"1f",x"fe"),
     6 => (x"48",x"d0",x"ff",x"1e"),
     7 => (x"71",x"78",x"c9",x"c8"),
     8 => (x"08",x"d4",x"ff",x"48"),
     9 => (x"1e",x"4f",x"26",x"78"),
    10 => (x"eb",x"49",x"4a",x"71"),
    11 => (x"48",x"d0",x"ff",x"87"),
    12 => (x"4f",x"26",x"78",x"c8"),
    13 => (x"71",x"1e",x"73",x"1e"),
    14 => (x"f0",x"f9",x"c2",x"4b"),
    15 => (x"87",x"c3",x"02",x"bf"),
    16 => (x"ff",x"87",x"eb",x"c2"),
    17 => (x"c9",x"c8",x"48",x"d0"),
    18 => (x"c0",x"49",x"73",x"78"),
    19 => (x"d4",x"ff",x"b1",x"e0"),
    20 => (x"c2",x"78",x"71",x"48"),
    21 => (x"c0",x"48",x"e4",x"f9"),
    22 => (x"02",x"66",x"c8",x"78"),
    23 => (x"ff",x"c3",x"87",x"c5"),
    24 => (x"c0",x"87",x"c2",x"49"),
    25 => (x"ec",x"f9",x"c2",x"49"),
    26 => (x"02",x"66",x"cc",x"59"),
    27 => (x"d5",x"c5",x"87",x"c6"),
    28 => (x"87",x"c4",x"4a",x"d5"),
    29 => (x"4a",x"ff",x"ff",x"cf"),
    30 => (x"5a",x"f0",x"f9",x"c2"),
    31 => (x"48",x"f0",x"f9",x"c2"),
    32 => (x"87",x"c4",x"78",x"c1"),
    33 => (x"4c",x"26",x"4d",x"26"),
    34 => (x"4f",x"26",x"4b",x"26"),
    35 => (x"5c",x"5b",x"5e",x"0e"),
    36 => (x"4a",x"71",x"0e",x"5d"),
    37 => (x"bf",x"ec",x"f9",x"c2"),
    38 => (x"02",x"9a",x"72",x"4c"),
    39 => (x"c8",x"49",x"87",x"cb"),
    40 => (x"ea",x"c0",x"c2",x"91"),
    41 => (x"c4",x"83",x"71",x"4b"),
    42 => (x"ea",x"c4",x"c2",x"87"),
    43 => (x"13",x"4d",x"c0",x"4b"),
    44 => (x"c2",x"99",x"74",x"49"),
    45 => (x"b9",x"bf",x"e8",x"f9"),
    46 => (x"71",x"48",x"d4",x"ff"),
    47 => (x"2c",x"b7",x"c1",x"78"),
    48 => (x"ad",x"b7",x"c8",x"85"),
    49 => (x"c2",x"87",x"e8",x"04"),
    50 => (x"48",x"bf",x"e4",x"f9"),
    51 => (x"f9",x"c2",x"80",x"c8"),
    52 => (x"ef",x"fe",x"58",x"e8"),
    53 => (x"1e",x"73",x"1e",x"87"),
    54 => (x"4a",x"13",x"4b",x"71"),
    55 => (x"87",x"cb",x"02",x"9a"),
    56 => (x"e7",x"fe",x"49",x"72"),
    57 => (x"9a",x"4a",x"13",x"87"),
    58 => (x"fe",x"87",x"f5",x"05"),
    59 => (x"c2",x"1e",x"87",x"da"),
    60 => (x"49",x"bf",x"e4",x"f9"),
    61 => (x"48",x"e4",x"f9",x"c2"),
    62 => (x"c4",x"78",x"a1",x"c1"),
    63 => (x"03",x"a9",x"b7",x"c0"),
    64 => (x"d4",x"ff",x"87",x"db"),
    65 => (x"e8",x"f9",x"c2",x"48"),
    66 => (x"f9",x"c2",x"78",x"bf"),
    67 => (x"c2",x"49",x"bf",x"e4"),
    68 => (x"c1",x"48",x"e4",x"f9"),
    69 => (x"c0",x"c4",x"78",x"a1"),
    70 => (x"e5",x"04",x"a9",x"b7"),
    71 => (x"48",x"d0",x"ff",x"87"),
    72 => (x"f9",x"c2",x"78",x"c8"),
    73 => (x"78",x"c0",x"48",x"f0"),
    74 => (x"00",x"00",x"4f",x"26"),
    75 => (x"00",x"00",x"00",x"00"),
    76 => (x"00",x"00",x"00",x"00"),
    77 => (x"00",x"5f",x"5f",x"00"),
    78 => (x"03",x"00",x"00",x"00"),
    79 => (x"03",x"03",x"00",x"03"),
    80 => (x"7f",x"14",x"00",x"00"),
    81 => (x"7f",x"7f",x"14",x"7f"),
    82 => (x"24",x"00",x"00",x"14"),
    83 => (x"3a",x"6b",x"6b",x"2e"),
    84 => (x"6a",x"4c",x"00",x"12"),
    85 => (x"56",x"6c",x"18",x"36"),
    86 => (x"7e",x"30",x"00",x"32"),
    87 => (x"3a",x"77",x"59",x"4f"),
    88 => (x"00",x"00",x"40",x"68"),
    89 => (x"00",x"03",x"07",x"04"),
    90 => (x"00",x"00",x"00",x"00"),
    91 => (x"41",x"63",x"3e",x"1c"),
    92 => (x"00",x"00",x"00",x"00"),
    93 => (x"1c",x"3e",x"63",x"41"),
    94 => (x"2a",x"08",x"00",x"00"),
    95 => (x"3e",x"1c",x"1c",x"3e"),
    96 => (x"08",x"00",x"08",x"2a"),
    97 => (x"08",x"3e",x"3e",x"08"),
    98 => (x"00",x"00",x"00",x"08"),
    99 => (x"00",x"60",x"e0",x"80"),
   100 => (x"08",x"00",x"00",x"00"),
   101 => (x"08",x"08",x"08",x"08"),
   102 => (x"00",x"00",x"00",x"08"),
   103 => (x"00",x"60",x"60",x"00"),
   104 => (x"60",x"40",x"00",x"00"),
   105 => (x"06",x"0c",x"18",x"30"),
   106 => (x"3e",x"00",x"01",x"03"),
   107 => (x"7f",x"4d",x"59",x"7f"),
   108 => (x"04",x"00",x"00",x"3e"),
   109 => (x"00",x"7f",x"7f",x"06"),
   110 => (x"42",x"00",x"00",x"00"),
   111 => (x"4f",x"59",x"71",x"63"),
   112 => (x"22",x"00",x"00",x"46"),
   113 => (x"7f",x"49",x"49",x"63"),
   114 => (x"1c",x"18",x"00",x"36"),
   115 => (x"7f",x"7f",x"13",x"16"),
   116 => (x"27",x"00",x"00",x"10"),
   117 => (x"7d",x"45",x"45",x"67"),
   118 => (x"3c",x"00",x"00",x"39"),
   119 => (x"79",x"49",x"4b",x"7e"),
   120 => (x"01",x"00",x"00",x"30"),
   121 => (x"0f",x"79",x"71",x"01"),
   122 => (x"36",x"00",x"00",x"07"),
   123 => (x"7f",x"49",x"49",x"7f"),
   124 => (x"06",x"00",x"00",x"36"),
   125 => (x"3f",x"69",x"49",x"4f"),
   126 => (x"00",x"00",x"00",x"1e"),
   127 => (x"00",x"66",x"66",x"00"),
   128 => (x"00",x"00",x"00",x"00"),
   129 => (x"00",x"66",x"e6",x"80"),
   130 => (x"08",x"00",x"00",x"00"),
   131 => (x"22",x"14",x"14",x"08"),
   132 => (x"14",x"00",x"00",x"22"),
   133 => (x"14",x"14",x"14",x"14"),
   134 => (x"22",x"00",x"00",x"14"),
   135 => (x"08",x"14",x"14",x"22"),
   136 => (x"02",x"00",x"00",x"08"),
   137 => (x"0f",x"59",x"51",x"03"),
   138 => (x"7f",x"3e",x"00",x"06"),
   139 => (x"1f",x"55",x"5d",x"41"),
   140 => (x"7e",x"00",x"00",x"1e"),
   141 => (x"7f",x"09",x"09",x"7f"),
   142 => (x"7f",x"00",x"00",x"7e"),
   143 => (x"7f",x"49",x"49",x"7f"),
   144 => (x"1c",x"00",x"00",x"36"),
   145 => (x"41",x"41",x"63",x"3e"),
   146 => (x"7f",x"00",x"00",x"41"),
   147 => (x"3e",x"63",x"41",x"7f"),
   148 => (x"7f",x"00",x"00",x"1c"),
   149 => (x"41",x"49",x"49",x"7f"),
   150 => (x"7f",x"00",x"00",x"41"),
   151 => (x"01",x"09",x"09",x"7f"),
   152 => (x"3e",x"00",x"00",x"01"),
   153 => (x"7b",x"49",x"41",x"7f"),
   154 => (x"7f",x"00",x"00",x"7a"),
   155 => (x"7f",x"08",x"08",x"7f"),
   156 => (x"00",x"00",x"00",x"7f"),
   157 => (x"41",x"7f",x"7f",x"41"),
   158 => (x"20",x"00",x"00",x"00"),
   159 => (x"7f",x"40",x"40",x"60"),
   160 => (x"7f",x"7f",x"00",x"3f"),
   161 => (x"63",x"36",x"1c",x"08"),
   162 => (x"7f",x"00",x"00",x"41"),
   163 => (x"40",x"40",x"40",x"7f"),
   164 => (x"7f",x"7f",x"00",x"40"),
   165 => (x"7f",x"06",x"0c",x"06"),
   166 => (x"7f",x"7f",x"00",x"7f"),
   167 => (x"7f",x"18",x"0c",x"06"),
   168 => (x"3e",x"00",x"00",x"7f"),
   169 => (x"7f",x"41",x"41",x"7f"),
   170 => (x"7f",x"00",x"00",x"3e"),
   171 => (x"0f",x"09",x"09",x"7f"),
   172 => (x"7f",x"3e",x"00",x"06"),
   173 => (x"7e",x"7f",x"61",x"41"),
   174 => (x"7f",x"00",x"00",x"40"),
   175 => (x"7f",x"19",x"09",x"7f"),
   176 => (x"26",x"00",x"00",x"66"),
   177 => (x"7b",x"59",x"4d",x"6f"),
   178 => (x"01",x"00",x"00",x"32"),
   179 => (x"01",x"7f",x"7f",x"01"),
   180 => (x"3f",x"00",x"00",x"01"),
   181 => (x"7f",x"40",x"40",x"7f"),
   182 => (x"0f",x"00",x"00",x"3f"),
   183 => (x"3f",x"70",x"70",x"3f"),
   184 => (x"7f",x"7f",x"00",x"0f"),
   185 => (x"7f",x"30",x"18",x"30"),
   186 => (x"63",x"41",x"00",x"7f"),
   187 => (x"36",x"1c",x"1c",x"36"),
   188 => (x"03",x"01",x"41",x"63"),
   189 => (x"06",x"7c",x"7c",x"06"),
   190 => (x"71",x"61",x"01",x"03"),
   191 => (x"43",x"47",x"4d",x"59"),
   192 => (x"00",x"00",x"00",x"41"),
   193 => (x"41",x"41",x"7f",x"7f"),
   194 => (x"03",x"01",x"00",x"00"),
   195 => (x"30",x"18",x"0c",x"06"),
   196 => (x"00",x"00",x"40",x"60"),
   197 => (x"7f",x"7f",x"41",x"41"),
   198 => (x"0c",x"08",x"00",x"00"),
   199 => (x"0c",x"06",x"03",x"06"),
   200 => (x"80",x"80",x"00",x"08"),
   201 => (x"80",x"80",x"80",x"80"),
   202 => (x"00",x"00",x"00",x"80"),
   203 => (x"04",x"07",x"03",x"00"),
   204 => (x"20",x"00",x"00",x"00"),
   205 => (x"7c",x"54",x"54",x"74"),
   206 => (x"7f",x"00",x"00",x"78"),
   207 => (x"7c",x"44",x"44",x"7f"),
   208 => (x"38",x"00",x"00",x"38"),
   209 => (x"44",x"44",x"44",x"7c"),
   210 => (x"38",x"00",x"00",x"00"),
   211 => (x"7f",x"44",x"44",x"7c"),
   212 => (x"38",x"00",x"00",x"7f"),
   213 => (x"5c",x"54",x"54",x"7c"),
   214 => (x"04",x"00",x"00",x"18"),
   215 => (x"05",x"05",x"7f",x"7e"),
   216 => (x"18",x"00",x"00",x"00"),
   217 => (x"fc",x"a4",x"a4",x"bc"),
   218 => (x"7f",x"00",x"00",x"7c"),
   219 => (x"7c",x"04",x"04",x"7f"),
   220 => (x"00",x"00",x"00",x"78"),
   221 => (x"40",x"7d",x"3d",x"00"),
   222 => (x"80",x"00",x"00",x"00"),
   223 => (x"7d",x"fd",x"80",x"80"),
   224 => (x"7f",x"00",x"00",x"00"),
   225 => (x"6c",x"38",x"10",x"7f"),
   226 => (x"00",x"00",x"00",x"44"),
   227 => (x"40",x"7f",x"3f",x"00"),
   228 => (x"7c",x"7c",x"00",x"00"),
   229 => (x"7c",x"0c",x"18",x"0c"),
   230 => (x"7c",x"00",x"00",x"78"),
   231 => (x"7c",x"04",x"04",x"7c"),
   232 => (x"38",x"00",x"00",x"78"),
   233 => (x"7c",x"44",x"44",x"7c"),
   234 => (x"fc",x"00",x"00",x"38"),
   235 => (x"3c",x"24",x"24",x"fc"),
   236 => (x"18",x"00",x"00",x"18"),
   237 => (x"fc",x"24",x"24",x"3c"),
   238 => (x"7c",x"00",x"00",x"fc"),
   239 => (x"0c",x"04",x"04",x"7c"),
   240 => (x"48",x"00",x"00",x"08"),
   241 => (x"74",x"54",x"54",x"5c"),
   242 => (x"04",x"00",x"00",x"20"),
   243 => (x"44",x"44",x"7f",x"3f"),
   244 => (x"3c",x"00",x"00",x"00"),
   245 => (x"7c",x"40",x"40",x"7c"),
   246 => (x"1c",x"00",x"00",x"7c"),
   247 => (x"3c",x"60",x"60",x"3c"),
   248 => (x"7c",x"3c",x"00",x"1c"),
   249 => (x"7c",x"60",x"30",x"60"),
   250 => (x"6c",x"44",x"00",x"3c"),
   251 => (x"6c",x"38",x"10",x"38"),
   252 => (x"1c",x"00",x"00",x"44"),
   253 => (x"3c",x"60",x"e0",x"bc"),
   254 => (x"44",x"00",x"00",x"1c"),
   255 => (x"4c",x"5c",x"74",x"64"),
   256 => (x"08",x"00",x"00",x"44"),
   257 => (x"41",x"77",x"3e",x"08"),
   258 => (x"00",x"00",x"00",x"41"),
   259 => (x"00",x"7f",x"7f",x"00"),
   260 => (x"41",x"00",x"00",x"00"),
   261 => (x"08",x"3e",x"77",x"41"),
   262 => (x"01",x"02",x"00",x"08"),
   263 => (x"02",x"02",x"03",x"01"),
   264 => (x"7f",x"7f",x"00",x"01"),
   265 => (x"7f",x"7f",x"7f",x"7f"),
   266 => (x"08",x"08",x"00",x"7f"),
   267 => (x"3e",x"3e",x"1c",x"1c"),
   268 => (x"7f",x"7f",x"7f",x"7f"),
   269 => (x"1c",x"1c",x"3e",x"3e"),
   270 => (x"10",x"00",x"08",x"08"),
   271 => (x"18",x"7c",x"7c",x"18"),
   272 => (x"10",x"00",x"00",x"10"),
   273 => (x"30",x"7c",x"7c",x"30"),
   274 => (x"30",x"10",x"00",x"10"),
   275 => (x"1e",x"78",x"60",x"60"),
   276 => (x"66",x"42",x"00",x"06"),
   277 => (x"66",x"3c",x"18",x"3c"),
   278 => (x"38",x"78",x"00",x"42"),
   279 => (x"6c",x"c6",x"c2",x"6a"),
   280 => (x"00",x"60",x"00",x"38"),
   281 => (x"00",x"00",x"60",x"00"),
   282 => (x"5e",x"0e",x"00",x"60"),
   283 => (x"0e",x"5d",x"5c",x"5b"),
   284 => (x"c2",x"4c",x"71",x"1e"),
   285 => (x"4d",x"bf",x"c1",x"fa"),
   286 => (x"1e",x"c0",x"4b",x"c0"),
   287 => (x"c7",x"02",x"ab",x"74"),
   288 => (x"48",x"a6",x"c4",x"87"),
   289 => (x"87",x"c5",x"78",x"c0"),
   290 => (x"c1",x"48",x"a6",x"c4"),
   291 => (x"1e",x"66",x"c4",x"78"),
   292 => (x"df",x"ee",x"49",x"73"),
   293 => (x"c0",x"86",x"c8",x"87"),
   294 => (x"ef",x"ef",x"49",x"e0"),
   295 => (x"4a",x"a5",x"c4",x"87"),
   296 => (x"f0",x"f0",x"49",x"6a"),
   297 => (x"87",x"c6",x"f1",x"87"),
   298 => (x"83",x"c1",x"85",x"cb"),
   299 => (x"04",x"ab",x"b7",x"c8"),
   300 => (x"26",x"87",x"c7",x"ff"),
   301 => (x"4c",x"26",x"4d",x"26"),
   302 => (x"4f",x"26",x"4b",x"26"),
   303 => (x"c2",x"4a",x"71",x"1e"),
   304 => (x"c2",x"5a",x"c5",x"fa"),
   305 => (x"c7",x"48",x"c5",x"fa"),
   306 => (x"dd",x"fe",x"49",x"78"),
   307 => (x"1e",x"4f",x"26",x"87"),
   308 => (x"4a",x"71",x"1e",x"73"),
   309 => (x"03",x"aa",x"b7",x"c0"),
   310 => (x"e0",x"c2",x"87",x"d3"),
   311 => (x"c4",x"05",x"bf",x"ef"),
   312 => (x"c2",x"4b",x"c1",x"87"),
   313 => (x"c2",x"4b",x"c0",x"87"),
   314 => (x"c4",x"5b",x"f3",x"e0"),
   315 => (x"f3",x"e0",x"c2",x"87"),
   316 => (x"ef",x"e0",x"c2",x"5a"),
   317 => (x"9a",x"c1",x"4a",x"bf"),
   318 => (x"49",x"a2",x"c0",x"c1"),
   319 => (x"fc",x"87",x"e8",x"ec"),
   320 => (x"ef",x"e0",x"c2",x"48"),
   321 => (x"ef",x"fe",x"78",x"bf"),
   322 => (x"4a",x"71",x"1e",x"87"),
   323 => (x"72",x"1e",x"66",x"c4"),
   324 => (x"dd",x"df",x"ff",x"49"),
   325 => (x"4f",x"26",x"26",x"87"),
   326 => (x"ef",x"e0",x"c2",x"1e"),
   327 => (x"dc",x"ff",x"49",x"bf"),
   328 => (x"f9",x"c2",x"87",x"cd"),
   329 => (x"bf",x"e8",x"48",x"f9"),
   330 => (x"f5",x"f9",x"c2",x"78"),
   331 => (x"78",x"bf",x"ec",x"48"),
   332 => (x"bf",x"f9",x"f9",x"c2"),
   333 => (x"ff",x"c3",x"49",x"4a"),
   334 => (x"2a",x"b7",x"c8",x"99"),
   335 => (x"b0",x"71",x"48",x"72"),
   336 => (x"58",x"c1",x"fa",x"c2"),
   337 => (x"5e",x"0e",x"4f",x"26"),
   338 => (x"0e",x"5d",x"5c",x"5b"),
   339 => (x"c7",x"ff",x"4b",x"71"),
   340 => (x"f4",x"f9",x"c2",x"87"),
   341 => (x"73",x"50",x"c0",x"48"),
   342 => (x"f2",x"db",x"ff",x"49"),
   343 => (x"4c",x"49",x"70",x"87"),
   344 => (x"ee",x"cb",x"9c",x"c2"),
   345 => (x"87",x"cf",x"cb",x"49"),
   346 => (x"c2",x"4d",x"49",x"70"),
   347 => (x"bf",x"97",x"f4",x"f9"),
   348 => (x"87",x"e4",x"c1",x"05"),
   349 => (x"c2",x"49",x"66",x"d0"),
   350 => (x"99",x"bf",x"fd",x"f9"),
   351 => (x"d4",x"87",x"d7",x"05"),
   352 => (x"f9",x"c2",x"49",x"66"),
   353 => (x"05",x"99",x"bf",x"f5"),
   354 => (x"49",x"73",x"87",x"cc"),
   355 => (x"87",x"ff",x"da",x"ff"),
   356 => (x"c1",x"02",x"98",x"70"),
   357 => (x"4c",x"c1",x"87",x"c2"),
   358 => (x"75",x"87",x"fd",x"fd"),
   359 => (x"87",x"e3",x"ca",x"49"),
   360 => (x"c6",x"02",x"98",x"70"),
   361 => (x"f4",x"f9",x"c2",x"87"),
   362 => (x"c2",x"50",x"c1",x"48"),
   363 => (x"bf",x"97",x"f4",x"f9"),
   364 => (x"87",x"e4",x"c0",x"05"),
   365 => (x"bf",x"fd",x"f9",x"c2"),
   366 => (x"99",x"66",x"d0",x"49"),
   367 => (x"87",x"d6",x"ff",x"05"),
   368 => (x"bf",x"f5",x"f9",x"c2"),
   369 => (x"99",x"66",x"d4",x"49"),
   370 => (x"87",x"ca",x"ff",x"05"),
   371 => (x"d9",x"ff",x"49",x"73"),
   372 => (x"98",x"70",x"87",x"fd"),
   373 => (x"87",x"fe",x"fe",x"05"),
   374 => (x"d7",x"fb",x"48",x"74"),
   375 => (x"5b",x"5e",x"0e",x"87"),
   376 => (x"f4",x"0e",x"5d",x"5c"),
   377 => (x"4c",x"4d",x"c0",x"86"),
   378 => (x"c4",x"7e",x"bf",x"ec"),
   379 => (x"fa",x"c2",x"48",x"a6"),
   380 => (x"c1",x"78",x"bf",x"c1"),
   381 => (x"c7",x"1e",x"c0",x"1e"),
   382 => (x"87",x"ca",x"fd",x"49"),
   383 => (x"98",x"70",x"86",x"c8"),
   384 => (x"ff",x"87",x"ce",x"02"),
   385 => (x"87",x"c7",x"fb",x"49"),
   386 => (x"ff",x"49",x"da",x"c1"),
   387 => (x"c1",x"87",x"c0",x"d9"),
   388 => (x"f4",x"f9",x"c2",x"4d"),
   389 => (x"c3",x"02",x"bf",x"97"),
   390 => (x"87",x"c0",x"c9",x"87"),
   391 => (x"bf",x"f9",x"f9",x"c2"),
   392 => (x"ef",x"e0",x"c2",x"4b"),
   393 => (x"eb",x"c0",x"05",x"bf"),
   394 => (x"49",x"fd",x"c3",x"87"),
   395 => (x"87",x"df",x"d8",x"ff"),
   396 => (x"ff",x"49",x"fa",x"c3"),
   397 => (x"73",x"87",x"d8",x"d8"),
   398 => (x"99",x"ff",x"c3",x"49"),
   399 => (x"49",x"c0",x"1e",x"71"),
   400 => (x"73",x"87",x"c6",x"fb"),
   401 => (x"29",x"b7",x"c8",x"49"),
   402 => (x"49",x"c1",x"1e",x"71"),
   403 => (x"c8",x"87",x"fa",x"fa"),
   404 => (x"87",x"c1",x"c6",x"86"),
   405 => (x"bf",x"fd",x"f9",x"c2"),
   406 => (x"dd",x"02",x"9b",x"4b"),
   407 => (x"eb",x"e0",x"c2",x"87"),
   408 => (x"de",x"c7",x"49",x"bf"),
   409 => (x"05",x"98",x"70",x"87"),
   410 => (x"4b",x"c0",x"87",x"c4"),
   411 => (x"e0",x"c2",x"87",x"d2"),
   412 => (x"87",x"c3",x"c7",x"49"),
   413 => (x"58",x"ef",x"e0",x"c2"),
   414 => (x"e0",x"c2",x"87",x"c6"),
   415 => (x"78",x"c0",x"48",x"eb"),
   416 => (x"99",x"c2",x"49",x"73"),
   417 => (x"c3",x"87",x"ce",x"05"),
   418 => (x"d7",x"ff",x"49",x"eb"),
   419 => (x"49",x"70",x"87",x"c1"),
   420 => (x"c2",x"02",x"99",x"c2"),
   421 => (x"73",x"4c",x"fb",x"87"),
   422 => (x"05",x"99",x"c1",x"49"),
   423 => (x"f4",x"c3",x"87",x"ce"),
   424 => (x"ea",x"d6",x"ff",x"49"),
   425 => (x"c2",x"49",x"70",x"87"),
   426 => (x"87",x"c2",x"02",x"99"),
   427 => (x"49",x"73",x"4c",x"fa"),
   428 => (x"ce",x"05",x"99",x"c8"),
   429 => (x"49",x"f5",x"c3",x"87"),
   430 => (x"87",x"d3",x"d6",x"ff"),
   431 => (x"99",x"c2",x"49",x"70"),
   432 => (x"c2",x"87",x"d5",x"02"),
   433 => (x"02",x"bf",x"c5",x"fa"),
   434 => (x"c1",x"48",x"87",x"ca"),
   435 => (x"c9",x"fa",x"c2",x"88"),
   436 => (x"87",x"c2",x"c0",x"58"),
   437 => (x"4d",x"c1",x"4c",x"ff"),
   438 => (x"99",x"c4",x"49",x"73"),
   439 => (x"c3",x"87",x"ce",x"05"),
   440 => (x"d5",x"ff",x"49",x"f2"),
   441 => (x"49",x"70",x"87",x"e9"),
   442 => (x"dc",x"02",x"99",x"c2"),
   443 => (x"c5",x"fa",x"c2",x"87"),
   444 => (x"c7",x"48",x"7e",x"bf"),
   445 => (x"c0",x"03",x"a8",x"b7"),
   446 => (x"48",x"6e",x"87",x"cb"),
   447 => (x"fa",x"c2",x"80",x"c1"),
   448 => (x"c2",x"c0",x"58",x"c9"),
   449 => (x"c1",x"4c",x"fe",x"87"),
   450 => (x"49",x"fd",x"c3",x"4d"),
   451 => (x"87",x"ff",x"d4",x"ff"),
   452 => (x"99",x"c2",x"49",x"70"),
   453 => (x"87",x"d5",x"c0",x"02"),
   454 => (x"bf",x"c5",x"fa",x"c2"),
   455 => (x"87",x"c9",x"c0",x"02"),
   456 => (x"48",x"c5",x"fa",x"c2"),
   457 => (x"c2",x"c0",x"78",x"c0"),
   458 => (x"c1",x"4c",x"fd",x"87"),
   459 => (x"49",x"fa",x"c3",x"4d"),
   460 => (x"87",x"db",x"d4",x"ff"),
   461 => (x"99",x"c2",x"49",x"70"),
   462 => (x"87",x"d9",x"c0",x"02"),
   463 => (x"bf",x"c5",x"fa",x"c2"),
   464 => (x"a8",x"b7",x"c7",x"48"),
   465 => (x"87",x"c9",x"c0",x"03"),
   466 => (x"48",x"c5",x"fa",x"c2"),
   467 => (x"c2",x"c0",x"78",x"c7"),
   468 => (x"c1",x"4c",x"fc",x"87"),
   469 => (x"ac",x"b7",x"c0",x"4d"),
   470 => (x"87",x"d1",x"c0",x"03"),
   471 => (x"c1",x"4a",x"66",x"c4"),
   472 => (x"02",x"6a",x"82",x"d8"),
   473 => (x"6a",x"87",x"c6",x"c0"),
   474 => (x"73",x"49",x"74",x"4b"),
   475 => (x"c3",x"1e",x"c0",x"0f"),
   476 => (x"da",x"c1",x"1e",x"f0"),
   477 => (x"87",x"ce",x"f7",x"49"),
   478 => (x"98",x"70",x"86",x"c8"),
   479 => (x"87",x"e2",x"c0",x"02"),
   480 => (x"c2",x"48",x"a6",x"c8"),
   481 => (x"78",x"bf",x"c5",x"fa"),
   482 => (x"cb",x"49",x"66",x"c8"),
   483 => (x"48",x"66",x"c4",x"91"),
   484 => (x"7e",x"70",x"80",x"71"),
   485 => (x"c0",x"02",x"bf",x"6e"),
   486 => (x"bf",x"6e",x"87",x"c8"),
   487 => (x"49",x"66",x"c8",x"4b"),
   488 => (x"9d",x"75",x"0f",x"73"),
   489 => (x"87",x"c8",x"c0",x"02"),
   490 => (x"bf",x"c5",x"fa",x"c2"),
   491 => (x"87",x"fa",x"f2",x"49"),
   492 => (x"bf",x"f3",x"e0",x"c2"),
   493 => (x"87",x"dd",x"c0",x"02"),
   494 => (x"87",x"c7",x"c2",x"49"),
   495 => (x"c0",x"02",x"98",x"70"),
   496 => (x"fa",x"c2",x"87",x"d3"),
   497 => (x"f2",x"49",x"bf",x"c5"),
   498 => (x"49",x"c0",x"87",x"e0"),
   499 => (x"c2",x"87",x"c0",x"f4"),
   500 => (x"c0",x"48",x"f3",x"e0"),
   501 => (x"f3",x"8e",x"f4",x"78"),
   502 => (x"5e",x"0e",x"87",x"da"),
   503 => (x"0e",x"5d",x"5c",x"5b"),
   504 => (x"c2",x"4c",x"71",x"1e"),
   505 => (x"49",x"bf",x"c1",x"fa"),
   506 => (x"4d",x"a1",x"cd",x"c1"),
   507 => (x"69",x"81",x"d1",x"c1"),
   508 => (x"02",x"9c",x"74",x"7e"),
   509 => (x"a5",x"c4",x"87",x"cf"),
   510 => (x"c2",x"7b",x"74",x"4b"),
   511 => (x"49",x"bf",x"c1",x"fa"),
   512 => (x"6e",x"87",x"f9",x"f2"),
   513 => (x"05",x"9c",x"74",x"7b"),
   514 => (x"4b",x"c0",x"87",x"c4"),
   515 => (x"4b",x"c1",x"87",x"c2"),
   516 => (x"fa",x"f2",x"49",x"73"),
   517 => (x"02",x"66",x"d4",x"87"),
   518 => (x"da",x"49",x"87",x"c7"),
   519 => (x"c2",x"4a",x"70",x"87"),
   520 => (x"c2",x"4a",x"c0",x"87"),
   521 => (x"26",x"5a",x"f7",x"e0"),
   522 => (x"00",x"87",x"c9",x"f2"),
   523 => (x"00",x"00",x"00",x"00"),
   524 => (x"00",x"00",x"00",x"00"),
   525 => (x"1e",x"00",x"00",x"00"),
   526 => (x"c8",x"ff",x"4a",x"71"),
   527 => (x"a1",x"72",x"49",x"bf"),
   528 => (x"1e",x"4f",x"26",x"48"),
   529 => (x"89",x"bf",x"c8",x"ff"),
   530 => (x"c0",x"c0",x"c0",x"fe"),
   531 => (x"01",x"a9",x"c0",x"c0"),
   532 => (x"4a",x"c0",x"87",x"c4"),
   533 => (x"4a",x"c1",x"87",x"c2"),
   534 => (x"4f",x"26",x"48",x"72"),
   535 => (x"ea",x"e2",x"c2",x"1e"),
   536 => (x"b9",x"c1",x"49",x"bf"),
   537 => (x"59",x"ee",x"e2",x"c2"),
   538 => (x"c3",x"48",x"d4",x"ff"),
   539 => (x"d0",x"ff",x"78",x"ff"),
   540 => (x"78",x"e1",x"c0",x"48"),
   541 => (x"c1",x"48",x"d4",x"ff"),
   542 => (x"71",x"31",x"c4",x"78"),
   543 => (x"48",x"d0",x"ff",x"78"),
   544 => (x"26",x"78",x"e0",x"c0"),
   545 => (x"e2",x"c2",x"1e",x"4f"),
   546 => (x"f4",x"c2",x"1e",x"de"),
   547 => (x"fd",x"fd",x"49",x"e8"),
   548 => (x"86",x"c4",x"87",x"df"),
   549 => (x"c3",x"02",x"98",x"70"),
   550 => (x"87",x"c0",x"ff",x"87"),
   551 => (x"35",x"31",x"4f",x"26"),
   552 => (x"20",x"5a",x"48",x"4b"),
   553 => (x"46",x"43",x"20",x"20"),
   554 => (x"00",x"00",x"00",x"47"),
   555 => (x"5e",x"0e",x"00",x"00"),
   556 => (x"0e",x"5d",x"5c",x"5b"),
   557 => (x"bf",x"f5",x"f9",x"c2"),
   558 => (x"d7",x"e4",x"c2",x"4a"),
   559 => (x"72",x"4c",x"49",x"bf"),
   560 => (x"ff",x"4d",x"71",x"bc"),
   561 => (x"c0",x"87",x"de",x"c6"),
   562 => (x"d0",x"49",x"74",x"4b"),
   563 => (x"e7",x"c0",x"02",x"99"),
   564 => (x"48",x"d0",x"ff",x"87"),
   565 => (x"ff",x"78",x"e1",x"c8"),
   566 => (x"78",x"c5",x"48",x"d4"),
   567 => (x"99",x"d0",x"49",x"75"),
   568 => (x"c3",x"87",x"c3",x"02"),
   569 => (x"e7",x"c2",x"78",x"f0"),
   570 => (x"81",x"73",x"49",x"c4"),
   571 => (x"d4",x"ff",x"48",x"11"),
   572 => (x"d0",x"ff",x"78",x"08"),
   573 => (x"78",x"e0",x"c0",x"48"),
   574 => (x"83",x"2d",x"2c",x"c1"),
   575 => (x"ff",x"04",x"ab",x"c8"),
   576 => (x"c5",x"ff",x"87",x"c7"),
   577 => (x"e4",x"c2",x"87",x"d7"),
   578 => (x"f9",x"c2",x"48",x"d7"),
   579 => (x"26",x"78",x"bf",x"f5"),
   580 => (x"26",x"4c",x"26",x"4d"),
   581 => (x"00",x"4f",x"26",x"4b"),
   582 => (x"1e",x"00",x"00",x"00"),
   583 => (x"4b",x"c0",x"1e",x"73"),
   584 => (x"48",x"cc",x"e7",x"c1"),
   585 => (x"1e",x"c8",x"50",x"de"),
   586 => (x"49",x"c9",x"fa",x"c2"),
   587 => (x"87",x"cc",x"d5",x"fe"),
   588 => (x"1e",x"72",x"86",x"c4"),
   589 => (x"48",x"cd",x"e6",x"c2"),
   590 => (x"49",x"d1",x"fa",x"c2"),
   591 => (x"20",x"4a",x"a1",x"c4"),
   592 => (x"05",x"aa",x"71",x"41"),
   593 => (x"4a",x"26",x"87",x"f9"),
   594 => (x"49",x"d1",x"e6",x"c2"),
   595 => (x"87",x"c2",x"f9",x"fd"),
   596 => (x"02",x"9a",x"4a",x"70"),
   597 => (x"fe",x"49",x"87",x"c5"),
   598 => (x"72",x"87",x"eb",x"c7"),
   599 => (x"dd",x"e6",x"c2",x"1e"),
   600 => (x"d1",x"fa",x"c2",x"48"),
   601 => (x"4a",x"a1",x"c4",x"49"),
   602 => (x"aa",x"71",x"41",x"20"),
   603 => (x"26",x"87",x"f9",x"05"),
   604 => (x"c9",x"fa",x"c2",x"4a"),
   605 => (x"dc",x"d9",x"fe",x"49"),
   606 => (x"05",x"98",x"70",x"87"),
   607 => (x"e6",x"c2",x"87",x"c4"),
   608 => (x"49",x"c0",x"4b",x"e1"),
   609 => (x"87",x"e0",x"c5",x"fe"),
   610 => (x"c6",x"fe",x"48",x"73"),
   611 => (x"20",x"20",x"20",x"87"),
   612 => (x"54",x"4f",x"4a",x"00"),
   613 => (x"20",x"4f",x"47",x"45"),
   614 => (x"20",x"20",x"20",x"20"),
   615 => (x"43",x"52",x"41",x"00"),
   616 => (x"43",x"52",x"41",x"00"),
   617 => (x"74",x"6f",x"6e",x"20"),
   618 => (x"75",x"6f",x"66",x"20"),
   619 => (x"20",x"2e",x"64",x"6e"),
   620 => (x"64",x"61",x"6f",x"4c"),
   621 => (x"43",x"52",x"41",x"20"),
   622 => (x"e0",x"f0",x"1e",x"00"),
   623 => (x"87",x"ee",x"fb",x"87"),
   624 => (x"4f",x"26",x"87",x"f8"),
   625 => (x"25",x"26",x"1e",x"16"),
   626 => (x"3e",x"3d",x"36",x"2e"),
		others => (others => x"00")
	);
	signal q1_local : word_t;

	-- Altera Quartus attributes
	attribute ramstyle: string;
	attribute ramstyle of ram: signal is "no_rw_check";

begin  -- rtl

	addr1 <= to_integer(unsigned(addr(ADDR_WIDTH-1 downto 0)));

	-- Reorganize the read data from the RAM to match the output
	q(7 downto 0) <= q1_local(3);
	q(15 downto 8) <= q1_local(2);
	q(23 downto 16) <= q1_local(1);
	q(31 downto 24) <= q1_local(0);

	process(clk)
	begin
		if(rising_edge(clk)) then 
			if(we = '1') then
				-- edit this code if using other than four bytes per word
				if (bytesel(3) = '1') then
					ram(addr1)(3) <= d(7 downto 0);
				end if;
				if (bytesel(2) = '1') then
					ram(addr1)(2) <= d(15 downto 8);
				end if;
				if (bytesel(1) = '1') then
					ram(addr1)(1) <= d(23 downto 16);
				end if;
				if (bytesel(0) = '1') then
					ram(addr1)(0) <= d(31 downto 24);
				end if;
			end if;
			q1_local <= ram(addr1);
		end if;
	end process;
  
end rtl;

