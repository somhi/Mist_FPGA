library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity controller_rom1 is
generic	(
	ADDR_WIDTH : integer := 8; -- ROM's address width (words, not bytes)
	COL_WIDTH  : integer := 8;  -- Column width (8bit -> byte)
	NB_COL     : integer := 4  -- Number of columns in memory
	);
port (
	clk : in std_logic;
	reset_n : in std_logic := '1';
	addr : in std_logic_vector(ADDR_WIDTH-1 downto 0);
	q : out std_logic_vector(31 downto 0);
	-- Allow writes - defaults supplied to simplify projects that don't need to write.
	d : in std_logic_vector(31 downto 0) := X"00000000";
	we : in std_logic := '0';
	bytesel : in std_logic_vector(3 downto 0) := "1111"
);
end entity;

architecture arch of controller_rom1 is

-- type word_t is std_logic_vector(31 downto 0);
type ram_type is array (0 to 2 ** ADDR_WIDTH - 1) of std_logic_vector(NB_COL * COL_WIDTH - 1 downto 0);

signal ram : ram_type :=
(

     0 => x"0487da01",
     1 => x"580e87dd",
     2 => x"0e5a595e",
     3 => x"00002927",
     4 => x"4a260f00",
     5 => x"48264926",
     6 => x"082680ff",
     7 => x"002d274f",
     8 => x"274f0000",
     9 => x"0000002a",
    10 => x"fd004f4f",
    11 => x"d8fac287",
    12 => x"86c0c54e",
    13 => x"49d8fac2",
    14 => x"48cce7c2",
    15 => x"4040c089",
    16 => x"89d04040",
    17 => x"c187f603",
    18 => x"0087e9e5",
    19 => x"1e87fc98",
    20 => x"1e731e72",
    21 => x"02114812",
    22 => x"c34b87ca",
    23 => x"739b98df",
    24 => x"87f00288",
    25 => x"4a264b26",
    26 => x"731e4f26",
    27 => x"c11e721e",
    28 => x"87ca048b",
    29 => x"02114812",
    30 => x"028887c4",
    31 => x"4a2687f1",
    32 => x"4f264b26",
    33 => x"731e741e",
    34 => x"c11e721e",
    35 => x"87d0048b",
    36 => x"02114812",
    37 => x"c34c87ca",
    38 => x"749c98df",
    39 => x"87eb0288",
    40 => x"4b264a26",
    41 => x"4f264c26",
    42 => x"8148731e",
    43 => x"c502a973",
    44 => x"05531287",
    45 => x"4f2687f6",
    46 => x"4a66c41e",
    47 => x"51124871",
    48 => x"2687fb05",
    49 => x"48731e4f",
    50 => x"05a97381",
    51 => x"87f95372",
    52 => x"711e4f26",
    53 => x"4966c44a",
    54 => x"c888c148",
    55 => x"997158a6",
    56 => x"ff87d602",
    57 => x"ffc348d4",
    58 => x"c4526878",
    59 => x"c1484966",
    60 => x"58a6c888",
    61 => x"ea059971",
    62 => x"1e4f2687",
    63 => x"d4ff1e73",
    64 => x"7bffc34b",
    65 => x"ffc34a6b",
    66 => x"c8496b7b",
    67 => x"c3b17232",
    68 => x"4a6b7bff",
    69 => x"b27131c8",
    70 => x"6b7bffc3",
    71 => x"7232c849",
    72 => x"c44871b1",
    73 => x"264d2687",
    74 => x"264b264c",
    75 => x"5b5e0e4f",
    76 => x"710e5d5c",
    77 => x"4cd4ff4a",
    78 => x"ffc34972",
    79 => x"c27c7199",
    80 => x"05bfcce7",
    81 => x"66d087c8",
    82 => x"d430c948",
    83 => x"66d058a6",
    84 => x"c329d849",
    85 => x"7c7199ff",
    86 => x"d04966d0",
    87 => x"99ffc329",
    88 => x"66d07c71",
    89 => x"c329c849",
    90 => x"7c7199ff",
    91 => x"c34966d0",
    92 => x"7c7199ff",
    93 => x"29d04972",
    94 => x"7199ffc3",
    95 => x"c94b6c7c",
    96 => x"c34dfff0",
    97 => x"d005abff",
    98 => x"7cffc387",
    99 => x"8dc14b6c",
   100 => x"c387c602",
   101 => x"f002abff",
   102 => x"fe487387",
   103 => x"c01e87c7",
   104 => x"48d4ff49",
   105 => x"c178ffc3",
   106 => x"b7c8c381",
   107 => x"87f104a9",
   108 => x"731e4f26",
   109 => x"c487e71e",
   110 => x"c04bdff8",
   111 => x"f0ffc01e",
   112 => x"fd49f7c1",
   113 => x"86c487e7",
   114 => x"c005a8c1",
   115 => x"d4ff87ea",
   116 => x"78ffc348",
   117 => x"c0c0c0c1",
   118 => x"c01ec0c0",
   119 => x"e9c1f0e1",
   120 => x"87c9fd49",
   121 => x"987086c4",
   122 => x"ff87ca05",
   123 => x"ffc348d4",
   124 => x"cb48c178",
   125 => x"87e6fe87",
   126 => x"fe058bc1",
   127 => x"48c087fd",
   128 => x"1e87e6fc",
   129 => x"d4ff1e73",
   130 => x"78ffc348",
   131 => x"1ec04bd3",
   132 => x"c1f0ffc0",
   133 => x"d4fc49c1",
   134 => x"7086c487",
   135 => x"87ca0598",
   136 => x"c348d4ff",
   137 => x"48c178ff",
   138 => x"f1fd87cb",
   139 => x"058bc187",
   140 => x"c087dbff",
   141 => x"87f1fb48",
   142 => x"5c5b5e0e",
   143 => x"4cd4ff0e",
   144 => x"c687dbfd",
   145 => x"e1c01eea",
   146 => x"49c8c1f0",
   147 => x"c487defb",
   148 => x"02a8c186",
   149 => x"eafe87c8",
   150 => x"c148c087",
   151 => x"dafa87e2",
   152 => x"cf497087",
   153 => x"c699ffff",
   154 => x"c802a9ea",
   155 => x"87d3fe87",
   156 => x"cbc148c0",
   157 => x"7cffc387",
   158 => x"fc4bf1c0",
   159 => x"987087f4",
   160 => x"87ebc002",
   161 => x"ffc01ec0",
   162 => x"49fac1f0",
   163 => x"c487defa",
   164 => x"05987086",
   165 => x"ffc387d9",
   166 => x"c3496c7c",
   167 => x"7c7c7cff",
   168 => x"99c0c17c",
   169 => x"c187c402",
   170 => x"c087d548",
   171 => x"c287d148",
   172 => x"87c405ab",
   173 => x"87c848c0",
   174 => x"fe058bc1",
   175 => x"48c087fd",
   176 => x"1e87e4f9",
   177 => x"e7c21e73",
   178 => x"78c148cc",
   179 => x"d0ff4bc7",
   180 => x"fb78c248",
   181 => x"d0ff87c8",
   182 => x"c078c348",
   183 => x"d0e5c01e",
   184 => x"f949c0c1",
   185 => x"86c487c7",
   186 => x"c105a8c1",
   187 => x"abc24b87",
   188 => x"c087c505",
   189 => x"87f9c048",
   190 => x"ff058bc1",
   191 => x"f7fc87d0",
   192 => x"d0e7c287",
   193 => x"05987058",
   194 => x"1ec187cd",
   195 => x"c1f0ffc0",
   196 => x"d8f849d0",
   197 => x"ff86c487",
   198 => x"ffc348d4",
   199 => x"87fcc278",
   200 => x"58d4e7c2",
   201 => x"c248d0ff",
   202 => x"48d4ff78",
   203 => x"c178ffc3",
   204 => x"87f5f748",
   205 => x"5c5b5e0e",
   206 => x"4b710e5d",
   207 => x"eec54cc0",
   208 => x"ff4adfcd",
   209 => x"ffc348d4",
   210 => x"c3496878",
   211 => x"c005a9fe",
   212 => x"4d7087fd",
   213 => x"cc029b73",
   214 => x"1e66d087",
   215 => x"f1f54973",
   216 => x"d686c487",
   217 => x"48d0ff87",
   218 => x"c378d1c4",
   219 => x"66d07dff",
   220 => x"d488c148",
   221 => x"987058a6",
   222 => x"ff87f005",
   223 => x"ffc348d4",
   224 => x"9b737878",
   225 => x"ff87c505",
   226 => x"78d048d0",
   227 => x"c14c4ac1",
   228 => x"eefe058a",
   229 => x"f6487487",
   230 => x"731e87cb",
   231 => x"c04a711e",
   232 => x"48d4ff4b",
   233 => x"ff78ffc3",
   234 => x"c3c448d0",
   235 => x"48d4ff78",
   236 => x"7278ffc3",
   237 => x"f0ffc01e",
   238 => x"f549d1c1",
   239 => x"86c487ef",
   240 => x"d2059870",
   241 => x"1ec0c887",
   242 => x"fd4966cc",
   243 => x"86c487e6",
   244 => x"d0ff4b70",
   245 => x"7378c248",
   246 => x"87cdf548",
   247 => x"5c5b5e0e",
   248 => x"1ec00e5d",
   249 => x"c1f0ffc0",
   250 => x"c0f549c9",
   251 => x"c21ed287",
   252 => x"fc49d4e7",
   253 => x"86c887fe",
   254 => x"84c14cc0",
   255 => x"04acb7d2",
   256 => x"e7c287f8",
   257 => x"49bf97d4",
   258 => x"c199c0c3",
   259 => x"c005a9c0",
   260 => x"e7c287e7",
   261 => x"49bf97db",
   262 => x"e7c231d0",
   263 => x"4abf97dc",
   264 => x"b17232c8",
   265 => x"97dde7c2",
   266 => x"71b14abf",
   267 => x"ffffcf4c",
   268 => x"84c19cff",
   269 => x"e7c134ca",
   270 => x"dde7c287",
   271 => x"c149bf97",
   272 => x"c299c631",
   273 => x"bf97dee7",
   274 => x"2ab7c74a",
   275 => x"e7c2b172",
   276 => x"4abf97d9",
   277 => x"c29dcf4d",
   278 => x"bf97dae7",
   279 => x"ca9ac34a",
   280 => x"dbe7c232",
   281 => x"c24bbf97",
   282 => x"c2b27333",
   283 => x"bf97dce7",
   284 => x"9bc0c34b",
   285 => x"732bb7c6",
   286 => x"c181c2b2",
   287 => x"70307148",
   288 => x"7548c149",
   289 => x"724d7030",
   290 => x"7184c14c",
   291 => x"b7c0c894",
   292 => x"87cc06ad",
   293 => x"2db734c1",
   294 => x"adb7c0c8",
   295 => x"87f4ff01",
   296 => x"c0f24874",
   297 => x"5b5e0e87",
   298 => x"f80e5d5c",
   299 => x"faefc286",
   300 => x"c278c048",
   301 => x"c01ef2e7",
   302 => x"87defb49",
   303 => x"987086c4",
   304 => x"c087c505",
   305 => x"87cec948",
   306 => x"7ec14dc0",
   307 => x"bfe2f5c0",
   308 => x"e8e8c249",
   309 => x"4bc8714a",
   310 => x"7087cfee",
   311 => x"87c20598",
   312 => x"f5c07ec0",
   313 => x"c249bfde",
   314 => x"714ac4e9",
   315 => x"f9ed4bc8",
   316 => x"05987087",
   317 => x"7ec087c2",
   318 => x"fdc0026e",
   319 => x"f8eec287",
   320 => x"efc24dbf",
   321 => x"7ebf9ff0",
   322 => x"ead6c548",
   323 => x"87c705a8",
   324 => x"bff8eec2",
   325 => x"6e87ce4d",
   326 => x"d5e9ca48",
   327 => x"87c502a8",
   328 => x"f1c748c0",
   329 => x"f2e7c287",
   330 => x"f949751e",
   331 => x"86c487ec",
   332 => x"c5059870",
   333 => x"c748c087",
   334 => x"f5c087dc",
   335 => x"c249bfde",
   336 => x"714ac4e9",
   337 => x"e1ec4bc8",
   338 => x"05987087",
   339 => x"efc287c8",
   340 => x"78c148fa",
   341 => x"f5c087da",
   342 => x"c249bfe2",
   343 => x"714ae8e8",
   344 => x"c5ec4bc8",
   345 => x"02987087",
   346 => x"c087c5c0",
   347 => x"87e6c648",
   348 => x"97f0efc2",
   349 => x"d5c149bf",
   350 => x"cdc005a9",
   351 => x"f1efc287",
   352 => x"c249bf97",
   353 => x"c002a9ea",
   354 => x"48c087c5",
   355 => x"c287c7c6",
   356 => x"bf97f2e7",
   357 => x"e9c3487e",
   358 => x"cec002a8",
   359 => x"c3486e87",
   360 => x"c002a8eb",
   361 => x"48c087c5",
   362 => x"c287ebc5",
   363 => x"bf97fde7",
   364 => x"c0059949",
   365 => x"e7c287cc",
   366 => x"49bf97fe",
   367 => x"c002a9c2",
   368 => x"48c087c5",
   369 => x"c287cfc5",
   370 => x"bf97ffe7",
   371 => x"f6efc248",
   372 => x"484c7058",
   373 => x"efc288c1",
   374 => x"e8c258fa",
   375 => x"49bf97c0",
   376 => x"e8c28175",
   377 => x"4abf97c1",
   378 => x"a17232c8",
   379 => x"c7f4c27e",
   380 => x"c2786e48",
   381 => x"bf97c2e8",
   382 => x"58a6c848",
   383 => x"bffaefc2",
   384 => x"87d4c202",
   385 => x"bfdef5c0",
   386 => x"c4e9c249",
   387 => x"4bc8714a",
   388 => x"7087d7e9",
   389 => x"c5c00298",
   390 => x"c348c087",
   391 => x"efc287f8",
   392 => x"c24cbff2",
   393 => x"c25cdbf4",
   394 => x"bf97d7e8",
   395 => x"c231c849",
   396 => x"bf97d6e8",
   397 => x"c249a14a",
   398 => x"bf97d8e8",
   399 => x"7232d04a",
   400 => x"e8c249a1",
   401 => x"4abf97d9",
   402 => x"a17232d8",
   403 => x"9166c449",
   404 => x"bfc7f4c2",
   405 => x"cff4c281",
   406 => x"dfe8c259",
   407 => x"c84abf97",
   408 => x"dee8c232",
   409 => x"a24bbf97",
   410 => x"e0e8c24a",
   411 => x"d04bbf97",
   412 => x"4aa27333",
   413 => x"97e1e8c2",
   414 => x"9bcf4bbf",
   415 => x"a27333d8",
   416 => x"d3f4c24a",
   417 => x"cff4c25a",
   418 => x"8ac24abf",
   419 => x"f4c29274",
   420 => x"a17248d3",
   421 => x"87cac178",
   422 => x"97c4e8c2",
   423 => x"31c849bf",
   424 => x"97c3e8c2",
   425 => x"49a14abf",
   426 => x"59c2f0c2",
   427 => x"bffeefc2",
   428 => x"c731c549",
   429 => x"29c981ff",
   430 => x"59dbf4c2",
   431 => x"97c9e8c2",
   432 => x"32c84abf",
   433 => x"97c8e8c2",
   434 => x"4aa24bbf",
   435 => x"6e9266c4",
   436 => x"d7f4c282",
   437 => x"cff4c25a",
   438 => x"c278c048",
   439 => x"7248cbf4",
   440 => x"f4c278a1",
   441 => x"f4c248db",
   442 => x"c278bfcf",
   443 => x"c248dff4",
   444 => x"78bfd3f4",
   445 => x"bffaefc2",
   446 => x"87c9c002",
   447 => x"30c44874",
   448 => x"c9c07e70",
   449 => x"d7f4c287",
   450 => x"30c448bf",
   451 => x"efc27e70",
   452 => x"786e48fe",
   453 => x"8ef848c1",
   454 => x"4c264d26",
   455 => x"4f264b26",
   456 => x"5c5b5e0e",
   457 => x"4a710e5d",
   458 => x"bffaefc2",
   459 => x"7287cb02",
   460 => x"722bc74b",
   461 => x"9cffc14c",
   462 => x"4b7287c9",
   463 => x"4c722bc8",
   464 => x"c29cffc3",
   465 => x"83bfc7f4",
   466 => x"bfdaf5c0",
   467 => x"87d902ab",
   468 => x"5bdef5c0",
   469 => x"1ef2e7c2",
   470 => x"fdf04973",
   471 => x"7086c487",
   472 => x"87c50598",
   473 => x"e6c048c0",
   474 => x"faefc287",
   475 => x"87d202bf",
   476 => x"91c44974",
   477 => x"81f2e7c2",
   478 => x"ffcf4d69",
   479 => x"9dffffff",
   480 => x"497487cb",
   481 => x"e7c291c2",
   482 => x"699f81f2",
   483 => x"fe48754d",
   484 => x"5e0e87c6",
   485 => x"0e5d5c5b",
   486 => x"c04d711e",
   487 => x"cf49c11e",
   488 => x"86c487dc",
   489 => x"029c4c70",
   490 => x"c287c0c1",
   491 => x"754ac2f0",
   492 => x"87dbe249",
   493 => x"c0029870",
   494 => x"4a7487f1",
   495 => x"4bcb4975",
   496 => x"7087c1e3",
   497 => x"e2c00298",
   498 => x"741ec087",
   499 => x"87c7029c",
   500 => x"c048a6c4",
   501 => x"c487c578",
   502 => x"78c148a6",
   503 => x"ce4966c4",
   504 => x"86c487dc",
   505 => x"059c4c70",
   506 => x"7487c0ff",
   507 => x"e7fc2648",
   508 => x"5b5e0e87",
   509 => x"1e0e5d5c",
   510 => x"059b4b71",
   511 => x"48c087c5",
   512 => x"c887e5c1",
   513 => x"7dc04da3",
   514 => x"c70266d4",
   515 => x"9766d487",
   516 => x"87c505bf",
   517 => x"cfc148c0",
   518 => x"4966d487",
   519 => x"7087f3fd",
   520 => x"c1029c4c",
   521 => x"a4dc87c0",
   522 => x"da7d6949",
   523 => x"a3c449a4",
   524 => x"7a699f4a",
   525 => x"bffaefc2",
   526 => x"d487d202",
   527 => x"699f49a4",
   528 => x"ffffc049",
   529 => x"d0487199",
   530 => x"c27e7030",
   531 => x"6e7ec087",
   532 => x"806a4849",
   533 => x"7bc07a70",
   534 => x"6a49a3cc",
   535 => x"49a3d079",
   536 => x"48c179c0",
   537 => x"48c087c2",
   538 => x"87ecfa26",
   539 => x"5c5b5e0e",
   540 => x"4c710e5d",
   541 => x"cac1029c",
   542 => x"49a4c887",
   543 => x"c2c10269",
   544 => x"4a66d087",
   545 => x"d482496c",
   546 => x"66d05aa6",
   547 => x"efc2b94d",
   548 => x"ff4abff6",
   549 => x"719972ba",
   550 => x"e4c00299",
   551 => x"4ba4c487",
   552 => x"fbf9496b",
   553 => x"c27b7087",
   554 => x"49bff2ef",
   555 => x"7c71816c",
   556 => x"efc2b975",
   557 => x"ff4abff6",
   558 => x"719972ba",
   559 => x"dcff0599",
   560 => x"f97c7587",
   561 => x"731e87d2",
   562 => x"9b4b711e",
   563 => x"c887c702",
   564 => x"056949a3",
   565 => x"48c087c5",
   566 => x"c287f7c0",
   567 => x"4abfcbf4",
   568 => x"6949a3c4",
   569 => x"c289c249",
   570 => x"91bff2ef",
   571 => x"c24aa271",
   572 => x"49bff6ef",
   573 => x"a271996b",
   574 => x"def5c04a",
   575 => x"1e66c85a",
   576 => x"d5ea4972",
   577 => x"7086c487",
   578 => x"87c40598",
   579 => x"87c248c0",
   580 => x"c7f848c1",
   581 => x"5b5e0e87",
   582 => x"1e0e5d5c",
   583 => x"66d44b71",
   584 => x"732cc94c",
   585 => x"cfc1029b",
   586 => x"49a3c887",
   587 => x"c7c10269",
   588 => x"4da3d087",
   589 => x"c27d66d4",
   590 => x"49bff6ef",
   591 => x"4a6bb9ff",
   592 => x"ac717e99",
   593 => x"c087cd03",
   594 => x"a3cc7d7b",
   595 => x"49a3c44a",
   596 => x"87c2796a",
   597 => x"9c748c72",
   598 => x"4987dd02",
   599 => x"fc49731e",
   600 => x"86c487ca",
   601 => x"c74966d4",
   602 => x"cb0299ff",
   603 => x"f2e7c287",
   604 => x"fd49731e",
   605 => x"86c487d0",
   606 => x"87dcf626",
   607 => x"5c5b5e0e",
   608 => x"86f00e5d",
   609 => x"c059a6d0",
   610 => x"cc4b66e4",
   611 => x"87ca0266",
   612 => x"7080c848",
   613 => x"05bf6e7e",
   614 => x"48c087c5",
   615 => x"cc87ecc3",
   616 => x"84d04c66",
   617 => x"a6c44973",
   618 => x"c4786c48",
   619 => x"80c48166",
   620 => x"c878bf6e",
   621 => x"c606a966",
   622 => x"66c44987",
   623 => x"c04b7189",
   624 => x"c401abb7",
   625 => x"c2c34887",
   626 => x"4866c487",
   627 => x"7098ffc7",
   628 => x"c1026e7e",
   629 => x"c0c887c9",
   630 => x"71896e49",
   631 => x"f2e7c24a",
   632 => x"73856e4d",
   633 => x"c106aab7",
   634 => x"49724a87",
   635 => x"8066c448",
   636 => x"8b727c70",
   637 => x"718ac149",
   638 => x"87d90299",
   639 => x"4866e0c0",
   640 => x"e0c05015",
   641 => x"80c14866",
   642 => x"58a6e4c0",
   643 => x"8ac14972",
   644 => x"e7059971",
   645 => x"d01ec187",
   646 => x"cff94966",
   647 => x"c086c487",
   648 => x"c106abb7",
   649 => x"e0c087e3",
   650 => x"ffc74d66",
   651 => x"c006abb7",
   652 => x"1e7587e2",
   653 => x"fa4966d0",
   654 => x"c0c887cc",
   655 => x"c8486c85",
   656 => x"7c7080c0",
   657 => x"c18bc0c8",
   658 => x"4966d41e",
   659 => x"c887ddf8",
   660 => x"87eec086",
   661 => x"1ef2e7c2",
   662 => x"f94966d0",
   663 => x"86c487e8",
   664 => x"4af2e7c2",
   665 => x"6c484973",
   666 => x"737c7080",
   667 => x"718bc149",
   668 => x"87ce0299",
   669 => x"c17d9712",
   670 => x"c1497385",
   671 => x"0599718b",
   672 => x"b7c087f2",
   673 => x"e1fe01ab",
   674 => x"f048c187",
   675 => x"87c8f28e",
   676 => x"5c5b5e0e",
   677 => x"4b710e5d",
   678 => x"87c7029b",
   679 => x"6d4da3c8",
   680 => x"ff87c505",
   681 => x"87fdc048",
   682 => x"6c4ca3d0",
   683 => x"99ffc749",
   684 => x"6c87d805",
   685 => x"c187c902",
   686 => x"f649731e",
   687 => x"86c487ee",
   688 => x"1ef2e7c2",
   689 => x"fdf74973",
   690 => x"6c86c487",
   691 => x"04aa6d4a",
   692 => x"48ff87c4",
   693 => x"a2c187cf",
   694 => x"c749727c",
   695 => x"e7c299ff",
   696 => x"699781f2",
   697 => x"87f0f048",
   698 => x"711e731e",
   699 => x"c0029b4b",
   700 => x"f4c287e4",
   701 => x"4a735bdf",
   702 => x"efc28ac2",
   703 => x"9249bff2",
   704 => x"bfcbf4c2",
   705 => x"c2807248",
   706 => x"7158e3f4",
   707 => x"c230c448",
   708 => x"c058c2f0",
   709 => x"f4c287ed",
   710 => x"f4c248db",
   711 => x"c278bfcf",
   712 => x"c248dff4",
   713 => x"78bfd3f4",
   714 => x"bffaefc2",
   715 => x"c287c902",
   716 => x"49bff2ef",
   717 => x"87c731c4",
   718 => x"bfd7f4c2",
   719 => x"c231c449",
   720 => x"ef59c2f0",
   721 => x"5e0e87d6",
   722 => x"710e5c5b",
   723 => x"724bc04a",
   724 => x"e1c0029a",
   725 => x"49a2da87",
   726 => x"c24b699f",
   727 => x"02bffaef",
   728 => x"a2d487cf",
   729 => x"49699f49",
   730 => x"ffffc04c",
   731 => x"c234d09c",
   732 => x"744cc087",
   733 => x"4973b349",
   734 => x"ee87edfd",
   735 => x"5e0e87dc",
   736 => x"0e5d5c5b",
   737 => x"4a7186f4",
   738 => x"9a727ec0",
   739 => x"c287d802",
   740 => x"c048eee7",
   741 => x"e6e7c278",
   742 => x"dff4c248",
   743 => x"e7c278bf",
   744 => x"f4c248ea",
   745 => x"c278bfdb",
   746 => x"c048cff0",
   747 => x"feefc250",
   748 => x"e7c249bf",
   749 => x"714abfee",
   750 => x"cac403aa",
   751 => x"cf497287",
   752 => x"eac00599",
   753 => x"daf5c087",
   754 => x"e6e7c248",
   755 => x"e7c278bf",
   756 => x"e7c21ef2",
   757 => x"c249bfe6",
   758 => x"c148e6e7",
   759 => x"ff7178a1",
   760 => x"c487f7de",
   761 => x"d6f5c086",
   762 => x"f2e7c248",
   763 => x"c087cc78",
   764 => x"48bfd6f5",
   765 => x"c080e0c0",
   766 => x"c258daf5",
   767 => x"48bfeee7",
   768 => x"e7c280c1",
   769 => x"562758f2",
   770 => x"bf00000d",
   771 => x"9d4dbf97",
   772 => x"87e3c202",
   773 => x"02ade5c3",
   774 => x"c087dcc2",
   775 => x"4bbfd6f5",
   776 => x"1149a3cb",
   777 => x"05accf4c",
   778 => x"7587d2c1",
   779 => x"c199df49",
   780 => x"c291cd89",
   781 => x"c181c2f0",
   782 => x"51124aa3",
   783 => x"124aa3c3",
   784 => x"4aa3c551",
   785 => x"a3c75112",
   786 => x"c951124a",
   787 => x"51124aa3",
   788 => x"124aa3ce",
   789 => x"4aa3d051",
   790 => x"a3d25112",
   791 => x"d451124a",
   792 => x"51124aa3",
   793 => x"124aa3d6",
   794 => x"4aa3d851",
   795 => x"a3dc5112",
   796 => x"de51124a",
   797 => x"51124aa3",
   798 => x"fac07ec1",
   799 => x"c8497487",
   800 => x"ebc00599",
   801 => x"d0497487",
   802 => x"87d10599",
   803 => x"c00266dc",
   804 => x"497387cb",
   805 => x"700f66dc",
   806 => x"d3c00298",
   807 => x"c0056e87",
   808 => x"f0c287c6",
   809 => x"50c048c2",
   810 => x"bfd6f5c0",
   811 => x"87e1c248",
   812 => x"48cff0c2",
   813 => x"c27e50c0",
   814 => x"49bffeef",
   815 => x"bfeee7c2",
   816 => x"04aa714a",
   817 => x"c287f6fb",
   818 => x"05bfdff4",
   819 => x"c287c8c0",
   820 => x"02bffaef",
   821 => x"c287f8c1",
   822 => x"49bfeae7",
   823 => x"7087c1e9",
   824 => x"eee7c249",
   825 => x"48a6c459",
   826 => x"bfeae7c2",
   827 => x"faefc278",
   828 => x"d8c002bf",
   829 => x"4966c487",
   830 => x"ffffffcf",
   831 => x"02a999f8",
   832 => x"c087c5c0",
   833 => x"87e1c04c",
   834 => x"dcc04cc1",
   835 => x"4966c487",
   836 => x"99f8ffcf",
   837 => x"c8c002a9",
   838 => x"48a6c887",
   839 => x"c5c078c0",
   840 => x"48a6c887",
   841 => x"66c878c1",
   842 => x"059c744c",
   843 => x"c487e0c0",
   844 => x"89c24966",
   845 => x"bff2efc2",
   846 => x"f4c2914a",
   847 => x"c24abfcb",
   848 => x"7248e6e7",
   849 => x"e7c278a1",
   850 => x"78c048ee",
   851 => x"c087def9",
   852 => x"e78ef448",
   853 => x"000087c2",
   854 => x"ffff0000",
   855 => x"0d66ffff",
   856 => x"0d6f0000",
   857 => x"41460000",
   858 => x"20323354",
   859 => x"46002020",
   860 => x"36315441",
   861 => x"00202020",
   862 => x"e4f4c21e",
   863 => x"a8dd48bf",
   864 => x"c187c905",
   865 => x"7087d8c2",
   866 => x"87c84a49",
   867 => x"c348d4ff",
   868 => x"4a6878ff",
   869 => x"4f264872",
   870 => x"e4f4c21e",
   871 => x"a8dd48bf",
   872 => x"c187c605",
   873 => x"d987e4c1",
   874 => x"48d4ff87",
   875 => x"ff78ffc3",
   876 => x"e1c048d0",
   877 => x"48d4ff78",
   878 => x"f4c278d4",
   879 => x"d4ff48e3",
   880 => x"4f2650bf",
   881 => x"48d0ff1e",
   882 => x"2678e0c0",
   883 => x"e7fe1e4f",
   884 => x"99497087",
   885 => x"c087c602",
   886 => x"f105a9fb",
   887 => x"26487187",
   888 => x"5b5e0e4f",
   889 => x"4b710e5c",
   890 => x"cbfe4cc0",
   891 => x"99497087",
   892 => x"87f9c002",
   893 => x"02a9ecc0",
   894 => x"c087f2c0",
   895 => x"c002a9fb",
   896 => x"66cc87eb",
   897 => x"c703acb7",
   898 => x"0266d087",
   899 => x"537187c2",
   900 => x"c2029971",
   901 => x"fd84c187",
   902 => x"497087de",
   903 => x"87cd0299",
   904 => x"02a9ecc0",
   905 => x"fbc087c7",
   906 => x"d5ff05a9",
   907 => x"0266d087",
   908 => x"97c087c3",
   909 => x"a9ecc07b",
   910 => x"7487c405",
   911 => x"7487c54a",
   912 => x"8a0ac04a",
   913 => x"87c24872",
   914 => x"4c264d26",
   915 => x"4f264b26",
   916 => x"87e4fc1e",
   917 => x"f0c04970",
   918 => x"ca04a9b7",
   919 => x"b7f9c087",
   920 => x"87c301a9",
   921 => x"c189f0c0",
   922 => x"04a9b7c1",
   923 => x"dac187ca",
   924 => x"c301a9b7",
   925 => x"89f7c087",
   926 => x"4f264871",
   927 => x"5c5b5e0e",
   928 => x"fc4c710e",
   929 => x"1ec187d2",
   930 => x"741e66d0",
   931 => x"87d1fd49",
   932 => x"4b7086c8",
   933 => x"c087edfc",
   934 => x"c203abb7",
   935 => x"cc8b0b87",
   936 => x"03abb766",
   937 => x"a37487cf",
   938 => x"c083c149",
   939 => x"66cc51e0",
   940 => x"f104abb7",
   941 => x"49a37487",
   942 => x"cdfe51c0",
   943 => x"5b5e0e87",
   944 => x"4a710e5c",
   945 => x"724cd4ff",
   946 => x"87e9c049",
   947 => x"029b4b70",
   948 => x"8bc187c2",
   949 => x"c548d0ff",
   950 => x"7cd5c178",
   951 => x"31c64973",
   952 => x"97cce7c1",
   953 => x"71484abf",
   954 => x"ff7c70b0",
   955 => x"78c448d0",
   956 => x"d5fd4873",
   957 => x"5b5e0e87",
   958 => x"f40e5d5c",
   959 => x"c44c7186",
   960 => x"78c048a6",
   961 => x"6e7ea4c8",
   962 => x"c149bf97",
   963 => x"dd05a9c1",
   964 => x"49a4c987",
   965 => x"c1496997",
   966 => x"d105a9d2",
   967 => x"49a4ca87",
   968 => x"c1496997",
   969 => x"c505a9c3",
   970 => x"c248df87",
   971 => x"e7f987e1",
   972 => x"c04bc087",
   973 => x"bf97d4ff",
   974 => x"04a9c049",
   975 => x"ccfa87cf",
   976 => x"c083c187",
   977 => x"bf97d4ff",
   978 => x"f106ab49",
   979 => x"d4ffc087",
   980 => x"cf02bf97",
   981 => x"87e0f887",
   982 => x"02994970",
   983 => x"ecc087c6",
   984 => x"87f105a9",
   985 => x"cff84bc0",
   986 => x"f84d7087",
   987 => x"a6cc87ca",
   988 => x"87c4f858",
   989 => x"83c14a70",
   990 => x"49bf976e",
   991 => x"87c702ad",
   992 => x"05adffc0",
   993 => x"c987eac0",
   994 => x"699749a4",
   995 => x"a966c849",
   996 => x"4887c702",
   997 => x"05a8ffc0",
   998 => x"a4ca87d7",
   999 => x"49699749",
  1000 => x"87c602aa",
  1001 => x"05aaffc0",
  1002 => x"a6c487c7",
  1003 => x"d378c148",
  1004 => x"adecc087",
  1005 => x"c087c602",
  1006 => x"c705adfb",
  1007 => x"c44bc087",
  1008 => x"78c148a6",
  1009 => x"fe0266c4",
  1010 => x"f7f787dc",
  1011 => x"f4487387",
  1012 => x"87f4f98e",
  1013 => x"5b5e0e00",
  1014 => x"1e0e5d5c",
  1015 => x"d4ff4d71",
  1016 => x"c21e754b",
  1017 => x"e049e8f4",
  1018 => x"86c487c7",
  1019 => x"c4029870",
  1020 => x"f4c287c8",
  1021 => x"754cbff0",
  1022 => x"87c1fb49",
  1023 => x"c005a8de",
  1024 => x"497587eb",
  1025 => x"87f5f5c0",
  1026 => x"db029870",
  1027 => x"ccf9c287",
  1028 => x"e1c01ebf",
  1029 => x"c4f3c049",
  1030 => x"c186c487",
  1031 => x"c048cce7",
  1032 => x"d8f9c250",
  1033 => x"87edfe49",
  1034 => x"cfc348c1",
  1035 => x"48d0ff87",
  1036 => x"d6c178c5",
  1037 => x"754ac07b",
  1038 => x"7b1149a2",
  1039 => x"b7cb82c1",
  1040 => x"87f304aa",
  1041 => x"ffc34acc",
  1042 => x"c082c17b",
  1043 => x"04aab7e0",
  1044 => x"d0ff87f4",
  1045 => x"c378c448",
  1046 => x"78c57bff",
  1047 => x"c17bd3c1",
  1048 => x"7478c47b",
  1049 => x"c0c2029c",
  1050 => x"f2e7c287",
  1051 => x"4dc0c87e",
  1052 => x"acb7c08c",
  1053 => x"c887c603",
  1054 => x"c04da4c0",
  1055 => x"adc0c84c",
  1056 => x"c287dc05",
  1057 => x"bf97e3f4",
  1058 => x"0299d049",
  1059 => x"1ec087d1",
  1060 => x"49e8f4c2",
  1061 => x"c487efe0",
  1062 => x"4a497086",
  1063 => x"c287eec0",
  1064 => x"c21ef2e7",
  1065 => x"e049e8f4",
  1066 => x"86c487dc",
  1067 => x"ff4a4970",
  1068 => x"c5c848d0",
  1069 => x"7bd4c178",
  1070 => x"7bbf976e",
  1071 => x"80c1486e",
  1072 => x"8dc17e70",
  1073 => x"87f0ff05",
  1074 => x"c448d0ff",
  1075 => x"059a7278",
  1076 => x"48c087c5",
  1077 => x"c187e5c0",
  1078 => x"e8f4c21e",
  1079 => x"cbdeff49",
  1080 => x"7486c487",
  1081 => x"c0fe059c",
  1082 => x"48d0ff87",
  1083 => x"d3c178c5",
  1084 => x"c47bc07b",
  1085 => x"c048c178",
  1086 => x"48c087c2",
  1087 => x"264d2626",
  1088 => x"264b264c",
  1089 => x"5b5e0e4f",
  1090 => x"1e0e5d5c",
  1091 => x"4cc04b71",
  1092 => x"c004ab4d",
  1093 => x"fbc087e8",
  1094 => x"9d751ef5",
  1095 => x"c087c402",
  1096 => x"c187c24a",
  1097 => x"e949724a",
  1098 => x"86c487d4",
  1099 => x"84c17e70",
  1100 => x"87c2056e",
  1101 => x"85c14c73",
  1102 => x"ff06ac73",
  1103 => x"486e87d8",
  1104 => x"87f9fe26",
  1105 => x"c44a711e",
  1106 => x"87c50566",
  1107 => x"c4fa4972",
  1108 => x"0e4f2687",
  1109 => x"5d5c5b5e",
  1110 => x"4c711e0e",
  1111 => x"c291de49",
  1112 => x"714dd0f5",
  1113 => x"026d9785",
  1114 => x"c287dcc1",
  1115 => x"4abffcf4",
  1116 => x"49728274",
  1117 => x"7087cefe",
  1118 => x"c0026e7e",
  1119 => x"f5c287f2",
  1120 => x"4a6e4bc4",
  1121 => x"fcfe49cb",
  1122 => x"4b7487de",
  1123 => x"e7c193cb",
  1124 => x"83c483dc",
  1125 => x"7bcbc7c1",
  1126 => x"cbc14974",
  1127 => x"7b7587cc",
  1128 => x"97cde7c1",
  1129 => x"c21e49bf",
  1130 => x"fe49c4f5",
  1131 => x"86c487d6",
  1132 => x"cac14974",
  1133 => x"49c087f4",
  1134 => x"87d3ccc1",
  1135 => x"48e4f4c2",
  1136 => x"49c178c0",
  1137 => x"2687c4dd",
  1138 => x"4c87f2fc",
  1139 => x"6964616f",
  1140 => x"2e2e676e",
  1141 => x"5e0e002e",
  1142 => x"710e5c5b",
  1143 => x"f4c24a4b",
  1144 => x"7282bffc",
  1145 => x"87ddfc49",
  1146 => x"029c4c70",
  1147 => x"e54987c4",
  1148 => x"f4c287d4",
  1149 => x"78c048fc",
  1150 => x"cedc49c1",
  1151 => x"87fffb87",
  1152 => x"5c5b5e0e",
  1153 => x"86f40e5d",
  1154 => x"4df2e7c2",
  1155 => x"a6c44cc0",
  1156 => x"c278c048",
  1157 => x"49bffcf4",
  1158 => x"c106a9c0",
  1159 => x"e7c287c1",
  1160 => x"029848f2",
  1161 => x"c087f8c0",
  1162 => x"c81ef5fb",
  1163 => x"87c70266",
  1164 => x"c048a6c4",
  1165 => x"c487c578",
  1166 => x"78c148a6",
  1167 => x"e44966c4",
  1168 => x"86c487fc",
  1169 => x"84c14d70",
  1170 => x"c14866c4",
  1171 => x"58a6c880",
  1172 => x"bffcf4c2",
  1173 => x"c603ac49",
  1174 => x"059d7587",
  1175 => x"c087c8ff",
  1176 => x"029d754c",
  1177 => x"c087e0c3",
  1178 => x"c81ef5fb",
  1179 => x"87c70266",
  1180 => x"c048a6cc",
  1181 => x"cc87c578",
  1182 => x"78c148a6",
  1183 => x"e34966cc",
  1184 => x"86c487fc",
  1185 => x"026e7e70",
  1186 => x"6e87e9c2",
  1187 => x"9781cb49",
  1188 => x"99d04969",
  1189 => x"87d6c102",
  1190 => x"4ad6c7c1",
  1191 => x"91cb4974",
  1192 => x"81dce7c1",
  1193 => x"81c87972",
  1194 => x"7451ffc3",
  1195 => x"c291de49",
  1196 => x"714dd0f5",
  1197 => x"97c1c285",
  1198 => x"49a5c17d",
  1199 => x"c251e0c0",
  1200 => x"bf97c2f0",
  1201 => x"c187d202",
  1202 => x"4ba5c284",
  1203 => x"4ac2f0c2",
  1204 => x"f7fe49db",
  1205 => x"dbc187d2",
  1206 => x"49a5cd87",
  1207 => x"84c151c0",
  1208 => x"6e4ba5c2",
  1209 => x"fe49cb4a",
  1210 => x"c187fdf6",
  1211 => x"c5c187c6",
  1212 => x"49744ad3",
  1213 => x"e7c191cb",
  1214 => x"797281dc",
  1215 => x"97c2f0c2",
  1216 => x"87d802bf",
  1217 => x"91de4974",
  1218 => x"f5c284c1",
  1219 => x"83714bd0",
  1220 => x"4ac2f0c2",
  1221 => x"f6fe49dd",
  1222 => x"87d887ce",
  1223 => x"93de4b74",
  1224 => x"83d0f5c2",
  1225 => x"c049a3cb",
  1226 => x"7384c151",
  1227 => x"49cb4a6e",
  1228 => x"87f4f5fe",
  1229 => x"c14866c4",
  1230 => x"58a6c880",
  1231 => x"c003acc7",
  1232 => x"056e87c5",
  1233 => x"7487e0fc",
  1234 => x"f68ef448",
  1235 => x"731e87ef",
  1236 => x"494b711e",
  1237 => x"e7c191cb",
  1238 => x"a1c881dc",
  1239 => x"cce7c14a",
  1240 => x"c9501248",
  1241 => x"ffc04aa1",
  1242 => x"501248d4",
  1243 => x"e7c181ca",
  1244 => x"501148cd",
  1245 => x"97cde7c1",
  1246 => x"c01e49bf",
  1247 => x"87c4f749",
  1248 => x"48e4f4c2",
  1249 => x"49c178de",
  1250 => x"2687c0d6",
  1251 => x"1e87f2f5",
  1252 => x"cb494a71",
  1253 => x"dce7c191",
  1254 => x"1181c881",
  1255 => x"e8f4c248",
  1256 => x"fcf4c258",
  1257 => x"c178c048",
  1258 => x"87dfd549",
  1259 => x"c01e4f26",
  1260 => x"dac4c149",
  1261 => x"1e4f2687",
  1262 => x"d2029971",
  1263 => x"f1e8c187",
  1264 => x"f750c048",
  1265 => x"cfcec180",
  1266 => x"d5e7c140",
  1267 => x"c187ce78",
  1268 => x"c148ede8",
  1269 => x"fc78cee7",
  1270 => x"eecec180",
  1271 => x"0e4f2678",
  1272 => x"0e5c5b5e",
  1273 => x"cb4a4c71",
  1274 => x"dce7c192",
  1275 => x"49a2c882",
  1276 => x"974ba2c9",
  1277 => x"971e4b6b",
  1278 => x"ca1e4969",
  1279 => x"c0491282",
  1280 => x"c087fae4",
  1281 => x"87c3d449",
  1282 => x"c1c14974",
  1283 => x"8ef887dc",
  1284 => x"1e87ecf3",
  1285 => x"4b711e73",
  1286 => x"87c3ff49",
  1287 => x"fefe4973",
  1288 => x"87ddf387",
  1289 => x"711e731e",
  1290 => x"4aa3c64b",
  1291 => x"c187db02",
  1292 => x"87d6028a",
  1293 => x"dac1028a",
  1294 => x"c0028a87",
  1295 => x"028a87fc",
  1296 => x"8a87e1c0",
  1297 => x"c187cb02",
  1298 => x"49c787db",
  1299 => x"c187c0fd",
  1300 => x"f4c287de",
  1301 => x"c102bffc",
  1302 => x"c14887cb",
  1303 => x"c0f5c288",
  1304 => x"87c1c158",
  1305 => x"bfc0f5c2",
  1306 => x"87f9c002",
  1307 => x"bffcf4c2",
  1308 => x"c280c148",
  1309 => x"c058c0f5",
  1310 => x"f4c287eb",
  1311 => x"c649bffc",
  1312 => x"c0f5c289",
  1313 => x"a9b7c059",
  1314 => x"c287da03",
  1315 => x"c048fcf4",
  1316 => x"c287d278",
  1317 => x"02bfc0f5",
  1318 => x"f4c287cb",
  1319 => x"c648bffc",
  1320 => x"c0f5c280",
  1321 => x"d149c058",
  1322 => x"497387e1",
  1323 => x"87fafec0",
  1324 => x"1e87cef1",
  1325 => x"4b711e73",
  1326 => x"48e4f4c2",
  1327 => x"49c078dd",
  1328 => x"7387c8d1",
  1329 => x"e1fec049",
  1330 => x"87f5f087",
  1331 => x"5c5b5e0e",
  1332 => x"cc4c710e",
  1333 => x"4b741e66",
  1334 => x"e7c193cb",
  1335 => x"a3c483dc",
  1336 => x"fe496a4a",
  1337 => x"c187d1ef",
  1338 => x"c87bcecd",
  1339 => x"66d449a3",
  1340 => x"49a3c951",
  1341 => x"ca5166d8",
  1342 => x"66dc49a3",
  1343 => x"feef2651",
  1344 => x"5b5e0e87",
  1345 => x"ff0e5d5c",
  1346 => x"a6d886cc",
  1347 => x"48a6c859",
  1348 => x"80c478c0",
  1349 => x"7866c8c1",
  1350 => x"78c180c4",
  1351 => x"48c0f5c2",
  1352 => x"f4c278c1",
  1353 => x"de48bfe4",
  1354 => x"87cb05a8",
  1355 => x"7087d1f3",
  1356 => x"59a6cc49",
  1357 => x"e187d0ce",
  1358 => x"d0e287de",
  1359 => x"87f8e087",
  1360 => x"66d44c70",
  1361 => x"87cac105",
  1362 => x"c11e1ec0",
  1363 => x"ffe8c11e",
  1364 => x"fd49c01e",
  1365 => x"86d087f6",
  1366 => x"02acfbc0",
  1367 => x"c4c187d9",
  1368 => x"82c44a66",
  1369 => x"81c7496a",
  1370 => x"1ec15174",
  1371 => x"496a1ed8",
  1372 => x"ece181c8",
  1373 => x"c186c887",
  1374 => x"c04866c8",
  1375 => x"87c701a8",
  1376 => x"c148a6c8",
  1377 => x"c187ce78",
  1378 => x"c14866c8",
  1379 => x"58a6d088",
  1380 => x"f8e087c3",
  1381 => x"48a6d887",
  1382 => x"9c7478c2",
  1383 => x"87e3cc02",
  1384 => x"c14866c8",
  1385 => x"03a866cc",
  1386 => x"c487d8cc",
  1387 => x"78c048a6",
  1388 => x"78c080d8",
  1389 => x"87c0dfff",
  1390 => x"66d44c70",
  1391 => x"05a8dd48",
  1392 => x"a6dc87c6",
  1393 => x"7866d448",
  1394 => x"05acd0c1",
  1395 => x"ff87ebc0",
  1396 => x"ff87e5de",
  1397 => x"7087e1de",
  1398 => x"acecc04c",
  1399 => x"ff87c605",
  1400 => x"7087eadf",
  1401 => x"acd0c14c",
  1402 => x"d087c805",
  1403 => x"80c14866",
  1404 => x"c158a6d4",
  1405 => x"ff02acd0",
  1406 => x"e0c087d5",
  1407 => x"66d448a6",
  1408 => x"4866dc78",
  1409 => x"a866e0c0",
  1410 => x"87c9ca05",
  1411 => x"48a6e4c0",
  1412 => x"80c478c0",
  1413 => x"4d7478c0",
  1414 => x"028dfbc0",
  1415 => x"c987cfc9",
  1416 => x"87db028d",
  1417 => x"c1028dc2",
  1418 => x"8dc987f7",
  1419 => x"87d2c402",
  1420 => x"c1028dc4",
  1421 => x"8dc187c2",
  1422 => x"87c6c402",
  1423 => x"c887e9c8",
  1424 => x"91cb4966",
  1425 => x"8166c4c1",
  1426 => x"6a4aa1c4",
  1427 => x"c11e717e",
  1428 => x"c448fee3",
  1429 => x"a1cc4966",
  1430 => x"7141204a",
  1431 => x"f8ff05aa",
  1432 => x"26511087",
  1433 => x"f3d2c149",
  1434 => x"e0ddff79",
  1435 => x"c04c7087",
  1436 => x"c148a6e8",
  1437 => x"87f6c778",
  1438 => x"c048a6c4",
  1439 => x"dbff78f0",
  1440 => x"4c7087f6",
  1441 => x"02acecc0",
  1442 => x"c887c3c0",
  1443 => x"ecc05ca6",
  1444 => x"87cd02ac",
  1445 => x"87e0dbff",
  1446 => x"ecc04c70",
  1447 => x"f3ff05ac",
  1448 => x"acecc087",
  1449 => x"87c4c002",
  1450 => x"87ccdbff",
  1451 => x"d41e66c4",
  1452 => x"c01e4966",
  1453 => x"1e4966e0",
  1454 => x"1effe8c1",
  1455 => x"f84966d8",
  1456 => x"1ec087ca",
  1457 => x"e0c01eca",
  1458 => x"91cb4966",
  1459 => x"8166dcc1",
  1460 => x"c448a6d8",
  1461 => x"66d878a1",
  1462 => x"dcff49bf",
  1463 => x"86d887c3",
  1464 => x"06a8b7c0",
  1465 => x"c187cbc1",
  1466 => x"c81ede1e",
  1467 => x"ff49bf66",
  1468 => x"c887eedb",
  1469 => x"48497086",
  1470 => x"c08808c0",
  1471 => x"c058a6ec",
  1472 => x"c006a8b7",
  1473 => x"e8c087ec",
  1474 => x"b7dd4866",
  1475 => x"e1c003a8",
  1476 => x"49bf6e87",
  1477 => x"8166e8c0",
  1478 => x"c051e0c0",
  1479 => x"c14966e8",
  1480 => x"81bf6e81",
  1481 => x"c051c1c2",
  1482 => x"c24966e8",
  1483 => x"81bf6e81",
  1484 => x"66d851c0",
  1485 => x"dc80c148",
  1486 => x"d04858a6",
  1487 => x"c478c180",
  1488 => x"dcff87ec",
  1489 => x"ecc087ca",
  1490 => x"dcff58a6",
  1491 => x"f0c087c2",
  1492 => x"ecc058a6",
  1493 => x"c9c005a8",
  1494 => x"c048a687",
  1495 => x"c07866e8",
  1496 => x"d8ff87c4",
  1497 => x"66c887d2",
  1498 => x"c191cb49",
  1499 => x"714866c4",
  1500 => x"58a6c880",
  1501 => x"c84a66c4",
  1502 => x"4966c482",
  1503 => x"e8c081ca",
  1504 => x"ecc05166",
  1505 => x"81c14966",
  1506 => x"8966e8c0",
  1507 => x"307148c1",
  1508 => x"89c14970",
  1509 => x"c27a9771",
  1510 => x"49bfecf8",
  1511 => x"2966e8c0",
  1512 => x"484a6a97",
  1513 => x"f4c09871",
  1514 => x"66c458a6",
  1515 => x"6981c449",
  1516 => x"66e0c07e",
  1517 => x"a866dc48",
  1518 => x"87c8c002",
  1519 => x"c048a6dc",
  1520 => x"87c5c078",
  1521 => x"c148a6dc",
  1522 => x"1e66dc78",
  1523 => x"c81ee0c0",
  1524 => x"d8ff4966",
  1525 => x"86c887cb",
  1526 => x"b7c04c70",
  1527 => x"d6c106ac",
  1528 => x"74486e87",
  1529 => x"c07e7080",
  1530 => x"897449e0",
  1531 => x"e3c14b6e",
  1532 => x"fe714afb",
  1533 => x"6e87f1e2",
  1534 => x"7080c248",
  1535 => x"66e4c07e",
  1536 => x"c080c148",
  1537 => x"c058a6e8",
  1538 => x"c14966f0",
  1539 => x"02a97081",
  1540 => x"c087c5c0",
  1541 => x"87c2c04d",
  1542 => x"1e754dc1",
  1543 => x"c049a4c2",
  1544 => x"887148e0",
  1545 => x"c81e4970",
  1546 => x"d6ff4966",
  1547 => x"86c887f3",
  1548 => x"01a8b7c0",
  1549 => x"c087c6ff",
  1550 => x"c00266e4",
  1551 => x"66c487d3",
  1552 => x"c081c949",
  1553 => x"c45166e4",
  1554 => x"cfc14866",
  1555 => x"cec078df",
  1556 => x"4966c487",
  1557 => x"51c281c9",
  1558 => x"c14866c4",
  1559 => x"c078d3d0",
  1560 => x"c148a6e8",
  1561 => x"87c6c078",
  1562 => x"87e1d5ff",
  1563 => x"e8c04c70",
  1564 => x"f5c00266",
  1565 => x"4866c887",
  1566 => x"04a866cc",
  1567 => x"c887cbc0",
  1568 => x"80c14866",
  1569 => x"c058a6cc",
  1570 => x"66cc87e0",
  1571 => x"d088c148",
  1572 => x"d5c058a6",
  1573 => x"acc6c187",
  1574 => x"87c8c005",
  1575 => x"c14866d8",
  1576 => x"58a6dc80",
  1577 => x"87e5d4ff",
  1578 => x"66d04c70",
  1579 => x"d480c148",
  1580 => x"9c7458a6",
  1581 => x"87cbc002",
  1582 => x"c14866c8",
  1583 => x"04a866cc",
  1584 => x"ff87e8f3",
  1585 => x"c887fdd3",
  1586 => x"a8c74866",
  1587 => x"87e5c003",
  1588 => x"48c0f5c2",
  1589 => x"66c878c0",
  1590 => x"c191cb49",
  1591 => x"c48166c4",
  1592 => x"4a6a4aa1",
  1593 => x"c87952c0",
  1594 => x"80c14866",
  1595 => x"c758a6cc",
  1596 => x"dbff04a8",
  1597 => x"8eccff87",
  1598 => x"3a87c2e0",
  1599 => x"49440020",
  1600 => x"77532050",
  1601 => x"68637469",
  1602 => x"1e007365",
  1603 => x"4b711e73",
  1604 => x"87c6029b",
  1605 => x"48fcf4c2",
  1606 => x"1ec778c0",
  1607 => x"bffcf4c2",
  1608 => x"e7c11e49",
  1609 => x"f4c21edc",
  1610 => x"ef49bfe4",
  1611 => x"86cc87d3",
  1612 => x"bfe4f4c2",
  1613 => x"87ffe949",
  1614 => x"c8029b73",
  1615 => x"dce7c187",
  1616 => x"f7edc049",
  1617 => x"f8deff87",
  1618 => x"d1c71e87",
  1619 => x"fe49c187",
  1620 => x"e5fe87f9",
  1621 => x"987087ed",
  1622 => x"fe87cd02",
  1623 => x"7087c6ed",
  1624 => x"87c40298",
  1625 => x"87c24ac1",
  1626 => x"9a724ac0",
  1627 => x"c087ce05",
  1628 => x"dee6c11e",
  1629 => x"e1f9c049",
  1630 => x"fe86c487",
  1631 => x"c4fcc087",
  1632 => x"c11ec087",
  1633 => x"c049e9e6",
  1634 => x"c087cff9",
  1635 => x"cafec01e",
  1636 => x"c0497087",
  1637 => x"c387c3f9",
  1638 => x"8ef887c3",
  1639 => x"44534f26",
  1640 => x"69616620",
  1641 => x"2e64656c",
  1642 => x"6f6f4200",
  1643 => x"676e6974",
  1644 => x"002e2e2e",
  1645 => x"fcf4c21e",
  1646 => x"c278c048",
  1647 => x"c048e4f4",
  1648 => x"87c5fe78",
  1649 => x"87f1ffc0",
  1650 => x"4f2648c0",
  1651 => x"20800000",
  1652 => x"74697845",
  1653 => x"42208000",
  1654 => x"006b6361",
  1655 => x"0000138f",
  1656 => x"00002d50",
  1657 => x"8f000000",
  1658 => x"6e000013",
  1659 => x"0000002d",
  1660 => x"138f0000",
  1661 => x"2d8c0000",
  1662 => x"00000000",
  1663 => x"00138f00",
  1664 => x"002daa00",
  1665 => x"00000000",
  1666 => x"0000138f",
  1667 => x"00002dc8",
  1668 => x"8f000000",
  1669 => x"e6000013",
  1670 => x"0000002d",
  1671 => x"138f0000",
  1672 => x"2e040000",
  1673 => x"00000000",
  1674 => x"00138f00",
  1675 => x"00000000",
  1676 => x"00000000",
  1677 => x"00001424",
  1678 => x"00000000",
  1679 => x"4c000000",
  1680 => x"2064616f",
  1681 => x"1e002e2a",
  1682 => x"c048f0fe",
  1683 => x"7909cd78",
  1684 => x"1e4f2609",
  1685 => x"bff0fe1e",
  1686 => x"2626487e",
  1687 => x"f0fe1e4f",
  1688 => x"2678c148",
  1689 => x"f0fe1e4f",
  1690 => x"2678c048",
  1691 => x"4a711e4f",
  1692 => x"265252c0",
  1693 => x"5b5e0e4f",
  1694 => x"f40e5d5c",
  1695 => x"974d7186",
  1696 => x"a5c17e6d",
  1697 => x"486c974c",
  1698 => x"6e58a6c8",
  1699 => x"a866c448",
  1700 => x"ff87c505",
  1701 => x"87e6c048",
  1702 => x"c287caff",
  1703 => x"6c9749a5",
  1704 => x"4ba3714b",
  1705 => x"974b6b97",
  1706 => x"486e7e6c",
  1707 => x"a6c880c1",
  1708 => x"cc98c758",
  1709 => x"977058a6",
  1710 => x"87e1fe7c",
  1711 => x"8ef44873",
  1712 => x"4c264d26",
  1713 => x"4f264b26",
  1714 => x"5c5b5e0e",
  1715 => x"7186f40e",
  1716 => x"4a66d84c",
  1717 => x"c29affc3",
  1718 => x"6c974ba4",
  1719 => x"49a17349",
  1720 => x"6c975172",
  1721 => x"c1486e7e",
  1722 => x"58a6c880",
  1723 => x"a6cc98c7",
  1724 => x"f4547058",
  1725 => x"87caff8e",
  1726 => x"e8fd1e1e",
  1727 => x"4abfe087",
  1728 => x"c0e0c049",
  1729 => x"87cb0299",
  1730 => x"f8c21e72",
  1731 => x"f7fe49e2",
  1732 => x"fc86c487",
  1733 => x"7e7087fd",
  1734 => x"2687c2fd",
  1735 => x"c21e4f26",
  1736 => x"fd49e2f8",
  1737 => x"ebc187c7",
  1738 => x"dafc49f8",
  1739 => x"87c8c487",
  1740 => x"ff1e4f26",
  1741 => x"e1c848d0",
  1742 => x"48d4ff78",
  1743 => x"66c478c5",
  1744 => x"c387c302",
  1745 => x"66c878e0",
  1746 => x"ff87c602",
  1747 => x"f0c348d4",
  1748 => x"48d4ff78",
  1749 => x"d0ff7871",
  1750 => x"78e1c848",
  1751 => x"2678e0c0",
  1752 => x"5b5e0e4f",
  1753 => x"4c710e5c",
  1754 => x"49e2f8c2",
  1755 => x"7087c6fc",
  1756 => x"aab7c04a",
  1757 => x"87e3c204",
  1758 => x"05aae0c3",
  1759 => x"f0c187c9",
  1760 => x"78c148eb",
  1761 => x"c387d4c2",
  1762 => x"c905aaf0",
  1763 => x"e7f0c187",
  1764 => x"c178c148",
  1765 => x"f0c187f5",
  1766 => x"c702bfeb",
  1767 => x"c24b7287",
  1768 => x"87c2b3c0",
  1769 => x"9c744b72",
  1770 => x"c187d105",
  1771 => x"1ebfe7f0",
  1772 => x"bfebf0c1",
  1773 => x"fd49721e",
  1774 => x"86c887f8",
  1775 => x"bfe7f0c1",
  1776 => x"87e0c002",
  1777 => x"b7c44973",
  1778 => x"f2c19129",
  1779 => x"4a7381c7",
  1780 => x"92c29acf",
  1781 => x"307248c1",
  1782 => x"baff4a70",
  1783 => x"98694872",
  1784 => x"87db7970",
  1785 => x"b7c44973",
  1786 => x"f2c19129",
  1787 => x"4a7381c7",
  1788 => x"92c29acf",
  1789 => x"307248c3",
  1790 => x"69484a70",
  1791 => x"c17970b0",
  1792 => x"c048ebf0",
  1793 => x"e7f0c178",
  1794 => x"c278c048",
  1795 => x"f949e2f8",
  1796 => x"4a7087e3",
  1797 => x"03aab7c0",
  1798 => x"c087ddfd",
  1799 => x"2687c248",
  1800 => x"264c264d",
  1801 => x"004f264b",
  1802 => x"00000000",
  1803 => x"1e000000",
  1804 => x"fc494a71",
  1805 => x"4f2687eb",
  1806 => x"724ac01e",
  1807 => x"c191c449",
  1808 => x"c081c7f2",
  1809 => x"d082c179",
  1810 => x"ee04aab7",
  1811 => x"0e4f2687",
  1812 => x"5d5c5b5e",
  1813 => x"f84d710e",
  1814 => x"4a7587cb",
  1815 => x"922ab7c4",
  1816 => x"82c7f2c1",
  1817 => x"9ccf4c75",
  1818 => x"496a94c2",
  1819 => x"c32b744b",
  1820 => x"7448c29b",
  1821 => x"ff4c7030",
  1822 => x"714874bc",
  1823 => x"f77a7098",
  1824 => x"487387db",
  1825 => x"0087d8fe",
  1826 => x"00000000",
  1827 => x"00000000",
  1828 => x"00000000",
  1829 => x"00000000",
  1830 => x"00000000",
  1831 => x"00000000",
  1832 => x"00000000",
  1833 => x"00000000",
  1834 => x"00000000",
  1835 => x"00000000",
  1836 => x"00000000",
  1837 => x"00000000",
  1838 => x"00000000",
  1839 => x"00000000",
  1840 => x"00000000",
  1841 => x"1e000000",
  1842 => x"c848d0ff",
  1843 => x"487178e1",
  1844 => x"7808d4ff",
  1845 => x"ff4866c4",
  1846 => x"267808d4",
  1847 => x"4a711e4f",
  1848 => x"1e4966c4",
  1849 => x"deff4972",
  1850 => x"48d0ff87",
  1851 => x"2678e0c0",
  1852 => x"731e4f26",
  1853 => x"c84b711e",
  1854 => x"731e4966",
  1855 => x"a2e0c14a",
  1856 => x"87d9ff49",
  1857 => x"2687c426",
  1858 => x"264c264d",
  1859 => x"1e4f264b",
  1860 => x"c34ad4ff",
  1861 => x"d0ff7aff",
  1862 => x"78e1c048",
  1863 => x"f8c27ade",
  1864 => x"497abfec",
  1865 => x"7028c848",
  1866 => x"d048717a",
  1867 => x"717a7028",
  1868 => x"7028d848",
  1869 => x"48d0ff7a",
  1870 => x"2678e0c0",
  1871 => x"5b5e0e4f",
  1872 => x"710e5d5c",
  1873 => x"ecf8c24c",
  1874 => x"744b4dbf",
  1875 => x"9b66d02b",
  1876 => x"66d483c1",
  1877 => x"87c204ab",
  1878 => x"4a744bc0",
  1879 => x"724966d0",
  1880 => x"75b9ff31",
  1881 => x"72487399",
  1882 => x"484a7030",
  1883 => x"f8c2b071",
  1884 => x"dafe58f0",
  1885 => x"264d2687",
  1886 => x"264b264c",
  1887 => x"5b5e0e4f",
  1888 => x"1e0e5d5c",
  1889 => x"f8c24c71",
  1890 => x"4ac04bf0",
  1891 => x"fe49f4c0",
  1892 => x"7487f2cc",
  1893 => x"f0f8c21e",
  1894 => x"d4e9fe49",
  1895 => x"7086c487",
  1896 => x"c0029949",
  1897 => x"1ec487ea",
  1898 => x"c21e4da6",
  1899 => x"fe49f0f8",
  1900 => x"c887c9ef",
  1901 => x"02987086",
  1902 => x"4a7587d6",
  1903 => x"49c6f8c1",
  1904 => x"cafe4bc4",
  1905 => x"987087e4",
  1906 => x"c087ca02",
  1907 => x"87edc048",
  1908 => x"e8c048c0",
  1909 => x"87f3c087",
  1910 => x"7087c4c1",
  1911 => x"87c80298",
  1912 => x"7087fcc0",
  1913 => x"87f80598",
  1914 => x"bfd0f9c2",
  1915 => x"c287cc02",
  1916 => x"c248ecf8",
  1917 => x"78bfd0f9",
  1918 => x"c187d4fc",
  1919 => x"4d262648",
  1920 => x"4b264c26",
  1921 => x"415b4f26",
  1922 => x"1e004352",
  1923 => x"f8c21ec0",
  1924 => x"ebfe49f0",
  1925 => x"f9c287ff",
  1926 => x"78c048c8",
  1927 => x"0e4f2626",
  1928 => x"5d5c5b5e",
  1929 => x"c486f40e",
  1930 => x"78c048a6",
  1931 => x"bfc8f9c2",
  1932 => x"a8b7c348",
  1933 => x"c287d103",
  1934 => x"48bfc8f9",
  1935 => x"f9c280c1",
  1936 => x"fbc058cc",
  1937 => x"87e2c648",
  1938 => x"49f0f8c2",
  1939 => x"87c0f1fe",
  1940 => x"f9c24c70",
  1941 => x"c34abfc8",
  1942 => x"87d8028a",
  1943 => x"c5028ac1",
  1944 => x"028a87cb",
  1945 => x"8a87f6c2",
  1946 => x"87cdc102",
  1947 => x"e2c3028a",
  1948 => x"87e1c587",
  1949 => x"4a754dc0",
  1950 => x"c0c292c4",
  1951 => x"f9c282c8",
  1952 => x"807548c4",
  1953 => x"976e7e70",
  1954 => x"4b494bbf",
  1955 => x"a3c1486e",
  1956 => x"11816a50",
  1957 => x"58a6cc48",
  1958 => x"c402ac70",
  1959 => x"c0486e87",
  1960 => x"0566c850",
  1961 => x"f9c287c7",
  1962 => x"a5c448c8",
  1963 => x"c485c178",
  1964 => x"ff04adb7",
  1965 => x"dcc487c0",
  1966 => x"d4f9c287",
  1967 => x"b7c848bf",
  1968 => x"87d101a8",
  1969 => x"cc02acca",
  1970 => x"02accd87",
  1971 => x"b7c087c7",
  1972 => x"f3c003ac",
  1973 => x"d4f9c287",
  1974 => x"b7c84bbf",
  1975 => x"87d203ab",
  1976 => x"49d8f9c2",
  1977 => x"e0c08173",
  1978 => x"c883c151",
  1979 => x"ff04abb7",
  1980 => x"f9c287ee",
  1981 => x"d2c148e0",
  1982 => x"50cfc150",
  1983 => x"c050cdc1",
  1984 => x"c380e450",
  1985 => x"87cdc378",
  1986 => x"bfd4f9c2",
  1987 => x"80c14849",
  1988 => x"58d8f9c2",
  1989 => x"81a0c448",
  1990 => x"f8c25174",
  1991 => x"b7f0c087",
  1992 => x"87da04ac",
  1993 => x"acb7f9c0",
  1994 => x"c287d301",
  1995 => x"49bfccf9",
  1996 => x"4a7491ca",
  1997 => x"c28af0c0",
  1998 => x"7248ccf9",
  1999 => x"acca78a1",
  2000 => x"87c6c002",
  2001 => x"c205accd",
  2002 => x"f9c287cb",
  2003 => x"78c348c8",
  2004 => x"c087c2c2",
  2005 => x"04acb7f0",
  2006 => x"f9c087db",
  2007 => x"c001acb7",
  2008 => x"f9c287d3",
  2009 => x"d049bfd0",
  2010 => x"c04a7491",
  2011 => x"f9c28af0",
  2012 => x"a17248d0",
  2013 => x"b7c1c178",
  2014 => x"dbc004ac",
  2015 => x"b7c6c187",
  2016 => x"d3c001ac",
  2017 => x"d0f9c287",
  2018 => x"91d049bf",
  2019 => x"f7c04a74",
  2020 => x"d0f9c28a",
  2021 => x"78a17248",
  2022 => x"c002acca",
  2023 => x"accd87c6",
  2024 => x"87f1c005",
  2025 => x"48c8f9c2",
  2026 => x"e8c078c3",
  2027 => x"ace2c087",
  2028 => x"87c9c005",
  2029 => x"c048a6c4",
  2030 => x"d8c078fb",
  2031 => x"02acca87",
  2032 => x"cd87c6c0",
  2033 => x"c9c005ac",
  2034 => x"c8f9c287",
  2035 => x"c078c348",
  2036 => x"a6c887c3",
  2037 => x"acb7c05c",
  2038 => x"87c4c003",
  2039 => x"87cac048",
  2040 => x"f90266c4",
  2041 => x"c34887c6",
  2042 => x"8ef499ff",
  2043 => x"4387cff8",
  2044 => x"3d464e4f",
  2045 => x"444f4d00",
  2046 => x"4d414e00",
  2047 => x"45440045",
  others => ( x"00000000")
);

-- Xilinx Vivado attributes
attribute ram_style: string;
attribute ram_style of ram: signal is "block";

signal q_local : std_logic_vector((NB_COL * COL_WIDTH)-1 downto 0);

signal wea : std_logic_vector(NB_COL - 1 downto 0);

begin

	output:
	for i in 0 to NB_COL - 1 generate
		q((i + 1) * COL_WIDTH - 1 downto i * COL_WIDTH) <= q_local((i+1) * COL_WIDTH - 1 downto i * COL_WIDTH);
	end generate;
    
    -- Generate write enable signals
    -- The Block ram generator doesn't like it when the compare is done in the if statement it self.
    wea <= bytesel when we = '1' else (others => '0');

    process(clk)
    begin
        if rising_edge(clk) then
            q_local <= ram(to_integer(unsigned(addr)));
            for i in 0 to NB_COL - 1 loop
                if (wea(NB_COL-i-1) = '1') then
                    ram(to_integer(unsigned(addr)))((i + 1) * COL_WIDTH - 1 downto i * COL_WIDTH) <= d((i + 1) * COL_WIDTH - 1 downto i * COL_WIDTH);
                end if;
            end loop;
        end if;
    end process;

end arch;
