library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity controller_rom is
generic	(
	ADDR_WIDTH : integer := 8; -- ROM's address width (words, not bytes)
	COL_WIDTH  : integer := 8;  -- Column width (8bit -> byte)
	NB_COL     : integer := 4  -- Number of columns in memory
	);
port (
	clk : in std_logic;
	reset_n : in std_logic := '1';
	addr : in std_logic_vector(ADDR_WIDTH-1 downto 0);
	q : out std_logic_vector(31 downto 0);
	-- Allow writes - defaults supplied to simplify projects that don't need to write.
	d : in std_logic_vector(31 downto 0) := X"00000000";
	we : in std_logic := '0';
	bytesel : in std_logic_vector(3 downto 0) := "1111"
);
end entity;

architecture arch of controller_rom is

-- type word_t is std_logic_vector(31 downto 0);
type ram_type is array (0 to 2 ** ADDR_WIDTH - 1) of std_logic_vector(NB_COL * COL_WIDTH - 1 downto 0);

signal ram : ram_type :=
(

     0 => x"0487da01",
     1 => x"580e87dd",
     2 => x"0e5a595e",
     3 => x"00002927",
     4 => x"4a260f00",
     5 => x"48264926",
     6 => x"082680ff",
     7 => x"002d274f",
     8 => x"274f0000",
     9 => x"0000002a",
    10 => x"fd004f4f",
    11 => x"c0f7c287",
    12 => x"86c0c84e",
    13 => x"49c0f7c2",
    14 => x"48c0e4c2",
    15 => x"4040c089",
    16 => x"89d04040",
    17 => x"c187f603",
    18 => x"0087e0e5",
    19 => x"1e87fc98",
    20 => x"1e731e72",
    21 => x"02114812",
    22 => x"c34b87ca",
    23 => x"739b98df",
    24 => x"87f00288",
    25 => x"4a264b26",
    26 => x"731e4f26",
    27 => x"c11e721e",
    28 => x"87ca048b",
    29 => x"02114812",
    30 => x"028887c4",
    31 => x"4a2687f1",
    32 => x"4f264b26",
    33 => x"731e741e",
    34 => x"c11e721e",
    35 => x"87d0048b",
    36 => x"02114812",
    37 => x"c34c87ca",
    38 => x"749c98df",
    39 => x"87eb0288",
    40 => x"4b264a26",
    41 => x"4f264c26",
    42 => x"8148731e",
    43 => x"c502a973",
    44 => x"05531287",
    45 => x"4f2687f6",
    46 => x"8148731e",
    47 => x"7205a973",
    48 => x"2687f953",
    49 => x"4a711e4f",
    50 => x"484966c4",
    51 => x"a6c888c1",
    52 => x"02997158",
    53 => x"d4ff87d6",
    54 => x"78ffc348",
    55 => x"66c45268",
    56 => x"88c14849",
    57 => x"7158a6c8",
    58 => x"87ea0599",
    59 => x"731e4f26",
    60 => x"4bd4ff1e",
    61 => x"6b7bffc3",
    62 => x"7bffc34a",
    63 => x"32c8496b",
    64 => x"ffc3b172",
    65 => x"c84a6b7b",
    66 => x"c3b27131",
    67 => x"496b7bff",
    68 => x"b17232c8",
    69 => x"87c44871",
    70 => x"4c264d26",
    71 => x"4f264b26",
    72 => x"5c5b5e0e",
    73 => x"4a710e5d",
    74 => x"724cd4ff",
    75 => x"99ffc349",
    76 => x"e4c27c71",
    77 => x"c805bfc0",
    78 => x"4866d087",
    79 => x"a6d430c9",
    80 => x"4966d058",
    81 => x"ffc329d8",
    82 => x"d07c7199",
    83 => x"29d04966",
    84 => x"7199ffc3",
    85 => x"4966d07c",
    86 => x"ffc329c8",
    87 => x"d07c7199",
    88 => x"ffc34966",
    89 => x"727c7199",
    90 => x"c329d049",
    91 => x"7c7199ff",
    92 => x"f0c94b6c",
    93 => x"ffc34dff",
    94 => x"87d005ab",
    95 => x"6c7cffc3",
    96 => x"028dc14b",
    97 => x"ffc387c6",
    98 => x"87f002ab",
    99 => x"c7fe4873",
   100 => x"49c01e87",
   101 => x"c348d4ff",
   102 => x"81c178ff",
   103 => x"a9b7c8c3",
   104 => x"2687f104",
   105 => x"1e731e4f",
   106 => x"f8c487e7",
   107 => x"1ec04bdf",
   108 => x"c1f0ffc0",
   109 => x"e7fd49f7",
   110 => x"c186c487",
   111 => x"eac005a8",
   112 => x"48d4ff87",
   113 => x"c178ffc3",
   114 => x"c0c0c0c0",
   115 => x"e1c01ec0",
   116 => x"49e9c1f0",
   117 => x"c487c9fd",
   118 => x"05987086",
   119 => x"d4ff87ca",
   120 => x"78ffc348",
   121 => x"87cb48c1",
   122 => x"c187e6fe",
   123 => x"fdfe058b",
   124 => x"fc48c087",
   125 => x"731e87e6",
   126 => x"48d4ff1e",
   127 => x"d378ffc3",
   128 => x"c01ec04b",
   129 => x"c1c1f0ff",
   130 => x"87d4fc49",
   131 => x"987086c4",
   132 => x"ff87ca05",
   133 => x"ffc348d4",
   134 => x"cb48c178",
   135 => x"87f1fd87",
   136 => x"ff058bc1",
   137 => x"48c087db",
   138 => x"0e87f1fb",
   139 => x"0e5c5b5e",
   140 => x"fd4cd4ff",
   141 => x"eac687db",
   142 => x"f0e1c01e",
   143 => x"fb49c8c1",
   144 => x"86c487de",
   145 => x"c802a8c1",
   146 => x"87eafe87",
   147 => x"e2c148c0",
   148 => x"87dafa87",
   149 => x"ffcf4970",
   150 => x"eac699ff",
   151 => x"87c802a9",
   152 => x"c087d3fe",
   153 => x"87cbc148",
   154 => x"c07cffc3",
   155 => x"f4fc4bf1",
   156 => x"02987087",
   157 => x"c087ebc0",
   158 => x"f0ffc01e",
   159 => x"fa49fac1",
   160 => x"86c487de",
   161 => x"d9059870",
   162 => x"7cffc387",
   163 => x"ffc3496c",
   164 => x"7c7c7c7c",
   165 => x"0299c0c1",
   166 => x"48c187c4",
   167 => x"48c087d5",
   168 => x"abc287d1",
   169 => x"c087c405",
   170 => x"c187c848",
   171 => x"fdfe058b",
   172 => x"f948c087",
   173 => x"731e87e4",
   174 => x"c0e4c21e",
   175 => x"c778c148",
   176 => x"48d0ff4b",
   177 => x"c8fb78c2",
   178 => x"48d0ff87",
   179 => x"1ec078c3",
   180 => x"c1d0e5c0",
   181 => x"c7f949c0",
   182 => x"c186c487",
   183 => x"87c105a8",
   184 => x"05abc24b",
   185 => x"48c087c5",
   186 => x"c187f9c0",
   187 => x"d0ff058b",
   188 => x"87f7fc87",
   189 => x"58c4e4c2",
   190 => x"cd059870",
   191 => x"c01ec187",
   192 => x"d0c1f0ff",
   193 => x"87d8f849",
   194 => x"d4ff86c4",
   195 => x"78ffc348",
   196 => x"c287fcc2",
   197 => x"ff58c8e4",
   198 => x"78c248d0",
   199 => x"c348d4ff",
   200 => x"48c178ff",
   201 => x"0e87f5f7",
   202 => x"5d5c5b5e",
   203 => x"c04b710e",
   204 => x"cdeec54c",
   205 => x"d4ff4adf",
   206 => x"78ffc348",
   207 => x"fec34968",
   208 => x"fdc005a9",
   209 => x"734d7087",
   210 => x"87cc029b",
   211 => x"731e66d0",
   212 => x"87f1f549",
   213 => x"87d686c4",
   214 => x"c448d0ff",
   215 => x"ffc378d1",
   216 => x"4866d07d",
   217 => x"a6d488c1",
   218 => x"05987058",
   219 => x"d4ff87f0",
   220 => x"78ffc348",
   221 => x"059b7378",
   222 => x"d0ff87c5",
   223 => x"c178d048",
   224 => x"8ac14c4a",
   225 => x"87eefe05",
   226 => x"cbf64874",
   227 => x"1e731e87",
   228 => x"4bc04a71",
   229 => x"c348d4ff",
   230 => x"d0ff78ff",
   231 => x"78c3c448",
   232 => x"c348d4ff",
   233 => x"1e7278ff",
   234 => x"c1f0ffc0",
   235 => x"eff549d1",
   236 => x"7086c487",
   237 => x"87d20598",
   238 => x"cc1ec0c8",
   239 => x"e6fd4966",
   240 => x"7086c487",
   241 => x"48d0ff4b",
   242 => x"487378c2",
   243 => x"0e87cdf5",
   244 => x"5d5c5b5e",
   245 => x"c01ec00e",
   246 => x"c9c1f0ff",
   247 => x"87c0f549",
   248 => x"e4c21ed2",
   249 => x"fefc49c8",
   250 => x"c086c887",
   251 => x"d284c14c",
   252 => x"f804acb7",
   253 => x"c8e4c287",
   254 => x"c349bf97",
   255 => x"c0c199c0",
   256 => x"e7c005a9",
   257 => x"cfe4c287",
   258 => x"d049bf97",
   259 => x"d0e4c231",
   260 => x"c84abf97",
   261 => x"c2b17232",
   262 => x"bf97d1e4",
   263 => x"4c71b14a",
   264 => x"ffffffcf",
   265 => x"ca84c19c",
   266 => x"87e7c134",
   267 => x"97d1e4c2",
   268 => x"31c149bf",
   269 => x"e4c299c6",
   270 => x"4abf97d2",
   271 => x"722ab7c7",
   272 => x"cde4c2b1",
   273 => x"4d4abf97",
   274 => x"e4c29dcf",
   275 => x"4abf97ce",
   276 => x"32ca9ac3",
   277 => x"97cfe4c2",
   278 => x"33c24bbf",
   279 => x"e4c2b273",
   280 => x"4bbf97d0",
   281 => x"c69bc0c3",
   282 => x"b2732bb7",
   283 => x"48c181c2",
   284 => x"49703071",
   285 => x"307548c1",
   286 => x"4c724d70",
   287 => x"947184c1",
   288 => x"adb7c0c8",
   289 => x"c187cc06",
   290 => x"c82db734",
   291 => x"01adb7c0",
   292 => x"7487f4ff",
   293 => x"87c0f248",
   294 => x"5c5b5e0e",
   295 => x"86f80e5d",
   296 => x"48eeecc2",
   297 => x"e4c278c0",
   298 => x"49c01ee6",
   299 => x"c487defb",
   300 => x"05987086",
   301 => x"48c087c5",
   302 => x"c087cec9",
   303 => x"c07ec14d",
   304 => x"49bfcff5",
   305 => x"4adce5c2",
   306 => x"ee4bc871",
   307 => x"987087dc",
   308 => x"c087c205",
   309 => x"cbf5c07e",
   310 => x"e5c249bf",
   311 => x"c8714af8",
   312 => x"87c6ee4b",
   313 => x"c2059870",
   314 => x"6e7ec087",
   315 => x"87fdc002",
   316 => x"bfecebc2",
   317 => x"e4ecc24d",
   318 => x"487ebf9f",
   319 => x"a8ead6c5",
   320 => x"c287c705",
   321 => x"4dbfeceb",
   322 => x"486e87ce",
   323 => x"a8d5e9ca",
   324 => x"c087c502",
   325 => x"87f1c748",
   326 => x"1ee6e4c2",
   327 => x"ecf94975",
   328 => x"7086c487",
   329 => x"87c50598",
   330 => x"dcc748c0",
   331 => x"cbf5c087",
   332 => x"e5c249bf",
   333 => x"c8714af8",
   334 => x"87eeec4b",
   335 => x"c8059870",
   336 => x"eeecc287",
   337 => x"da78c148",
   338 => x"cff5c087",
   339 => x"e5c249bf",
   340 => x"c8714adc",
   341 => x"87d2ec4b",
   342 => x"c0029870",
   343 => x"48c087c5",
   344 => x"c287e6c6",
   345 => x"bf97e4ec",
   346 => x"a9d5c149",
   347 => x"87cdc005",
   348 => x"97e5ecc2",
   349 => x"eac249bf",
   350 => x"c5c002a9",
   351 => x"c648c087",
   352 => x"e4c287c7",
   353 => x"7ebf97e6",
   354 => x"a8e9c348",
   355 => x"87cec002",
   356 => x"ebc3486e",
   357 => x"c5c002a8",
   358 => x"c548c087",
   359 => x"e4c287eb",
   360 => x"49bf97f1",
   361 => x"ccc00599",
   362 => x"f2e4c287",
   363 => x"c249bf97",
   364 => x"c5c002a9",
   365 => x"c548c087",
   366 => x"e4c287cf",
   367 => x"48bf97f3",
   368 => x"58eaecc2",
   369 => x"c1484c70",
   370 => x"eeecc288",
   371 => x"f4e4c258",
   372 => x"7549bf97",
   373 => x"f5e4c281",
   374 => x"c84abf97",
   375 => x"7ea17232",
   376 => x"48fbf0c2",
   377 => x"e4c2786e",
   378 => x"48bf97f6",
   379 => x"c258a6c8",
   380 => x"02bfeeec",
   381 => x"c087d4c2",
   382 => x"49bfcbf5",
   383 => x"4af8e5c2",
   384 => x"e94bc871",
   385 => x"987087e4",
   386 => x"87c5c002",
   387 => x"f8c348c0",
   388 => x"e6ecc287",
   389 => x"f1c24cbf",
   390 => x"e5c25ccf",
   391 => x"49bf97cb",
   392 => x"e5c231c8",
   393 => x"4abf97ca",
   394 => x"e5c249a1",
   395 => x"4abf97cc",
   396 => x"a17232d0",
   397 => x"cde5c249",
   398 => x"d84abf97",
   399 => x"49a17232",
   400 => x"c29166c4",
   401 => x"81bffbf0",
   402 => x"59c3f1c2",
   403 => x"97d3e5c2",
   404 => x"32c84abf",
   405 => x"97d2e5c2",
   406 => x"4aa24bbf",
   407 => x"97d4e5c2",
   408 => x"33d04bbf",
   409 => x"c24aa273",
   410 => x"bf97d5e5",
   411 => x"d89bcf4b",
   412 => x"4aa27333",
   413 => x"5ac7f1c2",
   414 => x"bfc3f1c2",
   415 => x"748ac24a",
   416 => x"c7f1c292",
   417 => x"78a17248",
   418 => x"c287cac1",
   419 => x"bf97f8e4",
   420 => x"c231c849",
   421 => x"bf97f7e4",
   422 => x"c249a14a",
   423 => x"c259f6ec",
   424 => x"49bff2ec",
   425 => x"ffc731c5",
   426 => x"c229c981",
   427 => x"c259cff1",
   428 => x"bf97fde4",
   429 => x"c232c84a",
   430 => x"bf97fce4",
   431 => x"c44aa24b",
   432 => x"826e9266",
   433 => x"5acbf1c2",
   434 => x"48c3f1c2",
   435 => x"f0c278c0",
   436 => x"a17248ff",
   437 => x"cff1c278",
   438 => x"c3f1c248",
   439 => x"f1c278bf",
   440 => x"f1c248d3",
   441 => x"c278bfc7",
   442 => x"02bfeeec",
   443 => x"7487c9c0",
   444 => x"7030c448",
   445 => x"87c9c07e",
   446 => x"bfcbf1c2",
   447 => x"7030c448",
   448 => x"f2ecc27e",
   449 => x"c1786e48",
   450 => x"268ef848",
   451 => x"264c264d",
   452 => x"0e4f264b",
   453 => x"5d5c5b5e",
   454 => x"c24a710e",
   455 => x"02bfeeec",
   456 => x"4b7287cb",
   457 => x"4c722bc7",
   458 => x"c99cffc1",
   459 => x"c84b7287",
   460 => x"c34c722b",
   461 => x"f0c29cff",
   462 => x"c083bffb",
   463 => x"abbfc7f5",
   464 => x"c087d902",
   465 => x"c25bcbf5",
   466 => x"731ee6e4",
   467 => x"87fdf049",
   468 => x"987086c4",
   469 => x"c087c505",
   470 => x"87e6c048",
   471 => x"bfeeecc2",
   472 => x"7487d202",
   473 => x"c291c449",
   474 => x"6981e6e4",
   475 => x"ffffcf4d",
   476 => x"cb9dffff",
   477 => x"c2497487",
   478 => x"e6e4c291",
   479 => x"4d699f81",
   480 => x"c6fe4875",
   481 => x"5b5e0e87",
   482 => x"f80e5d5c",
   483 => x"9c4c7186",
   484 => x"c087c505",
   485 => x"87c1c348",
   486 => x"6e7ea4c8",
   487 => x"d878c048",
   488 => x"87c70266",
   489 => x"bf9766d8",
   490 => x"c087c505",
   491 => x"87e9c248",
   492 => x"49c11ec0",
   493 => x"c487f4ce",
   494 => x"9d4d7086",
   495 => x"87c2c102",
   496 => x"4af6ecc2",
   497 => x"e24966d8",
   498 => x"987087c5",
   499 => x"87f2c002",
   500 => x"66d84a75",
   501 => x"e24bcb49",
   502 => x"987087ea",
   503 => x"87e2c002",
   504 => x"9d751ec0",
   505 => x"c887c702",
   506 => x"78c048a6",
   507 => x"a6c887c5",
   508 => x"c878c148",
   509 => x"f2cd4966",
   510 => x"7086c487",
   511 => x"fe059d4d",
   512 => x"9d7587fe",
   513 => x"87cfc102",
   514 => x"6e49a5dc",
   515 => x"da786948",
   516 => x"a6c449a5",
   517 => x"78a4c448",
   518 => x"c448699f",
   519 => x"c2780866",
   520 => x"02bfeeec",
   521 => x"a5d487d2",
   522 => x"49699f49",
   523 => x"99ffffc0",
   524 => x"30d04871",
   525 => x"87c27e70",
   526 => x"496e7ec0",
   527 => x"bf66c448",
   528 => x"0866c480",
   529 => x"cc7cc078",
   530 => x"66c449a4",
   531 => x"a4d079bf",
   532 => x"c179c049",
   533 => x"c087c248",
   534 => x"fa8ef848",
   535 => x"5e0e87ed",
   536 => x"0e5d5c5b",
   537 => x"029c4c71",
   538 => x"c887cac1",
   539 => x"026949a4",
   540 => x"d087c2c1",
   541 => x"496c4a66",
   542 => x"5aa6d482",
   543 => x"b94d66d0",
   544 => x"bfeaecc2",
   545 => x"72baff4a",
   546 => x"02997199",
   547 => x"c487e4c0",
   548 => x"496b4ba4",
   549 => x"7087fcf9",
   550 => x"e6ecc27b",
   551 => x"816c49bf",
   552 => x"b9757c71",
   553 => x"bfeaecc2",
   554 => x"72baff4a",
   555 => x"05997199",
   556 => x"7587dcff",
   557 => x"87d3f97c",
   558 => x"711e731e",
   559 => x"c7029b4b",
   560 => x"49a3c887",
   561 => x"87c50569",
   562 => x"f7c048c0",
   563 => x"fff0c287",
   564 => x"a3c44abf",
   565 => x"c2496949",
   566 => x"e6ecc289",
   567 => x"a27191bf",
   568 => x"eaecc24a",
   569 => x"996b49bf",
   570 => x"c04aa271",
   571 => x"c85acbf5",
   572 => x"49721e66",
   573 => x"c487d6ea",
   574 => x"05987086",
   575 => x"48c087c4",
   576 => x"48c187c2",
   577 => x"0e87c8f8",
   578 => x"5d5c5b5e",
   579 => x"4b711e0e",
   580 => x"734d66d4",
   581 => x"ccc1029b",
   582 => x"49a3c887",
   583 => x"c4c10269",
   584 => x"4ca3d087",
   585 => x"bfeaecc2",
   586 => x"6cb9ff49",
   587 => x"d47e994a",
   588 => x"cd06a966",
   589 => x"7c7bc087",
   590 => x"c44aa3cc",
   591 => x"796a49a3",
   592 => x"497287ca",
   593 => x"d499c0f8",
   594 => x"8d714d66",
   595 => x"29c94975",
   596 => x"49731e71",
   597 => x"c287c7fc",
   598 => x"731ee6e4",
   599 => x"87d8fd49",
   600 => x"66d486c8",
   601 => x"e2f6267c",
   602 => x"5b5e0e87",
   603 => x"f00e5d5c",
   604 => x"59a6d086",
   605 => x"4b66e4c0",
   606 => x"ca0266cc",
   607 => x"80c84887",
   608 => x"bf6e7e70",
   609 => x"c087c505",
   610 => x"87ecc348",
   611 => x"d04c66cc",
   612 => x"c4497384",
   613 => x"786c48a6",
   614 => x"c48166c4",
   615 => x"78bf6e80",
   616 => x"06a966c8",
   617 => x"c44987c6",
   618 => x"4b718966",
   619 => x"01abb7c0",
   620 => x"c34887c4",
   621 => x"66c487c2",
   622 => x"98ffc748",
   623 => x"026e7e70",
   624 => x"c887c9c1",
   625 => x"896e49c0",
   626 => x"e4c24a71",
   627 => x"856e4de6",
   628 => x"06aab773",
   629 => x"724a87c1",
   630 => x"66c44849",
   631 => x"727c7080",
   632 => x"8ac1498b",
   633 => x"d9029971",
   634 => x"66e0c087",
   635 => x"c0501548",
   636 => x"c14866e0",
   637 => x"a6e4c080",
   638 => x"c1497258",
   639 => x"0599718a",
   640 => x"1ec187e7",
   641 => x"f94966d0",
   642 => x"86c487d4",
   643 => x"06abb7c0",
   644 => x"c087e3c1",
   645 => x"c74d66e0",
   646 => x"06abb7ff",
   647 => x"7587e2c0",
   648 => x"4966d01e",
   649 => x"c887d1fa",
   650 => x"486c85c0",
   651 => x"7080c0c8",
   652 => x"8bc0c87c",
   653 => x"66d41ec1",
   654 => x"87e2f849",
   655 => x"eec086c8",
   656 => x"e6e4c287",
   657 => x"4966d01e",
   658 => x"c487edf9",
   659 => x"e6e4c286",
   660 => x"4849734a",
   661 => x"7c70806c",
   662 => x"8bc14973",
   663 => x"ce029971",
   664 => x"7d971287",
   665 => x"497385c1",
   666 => x"99718bc1",
   667 => x"c087f205",
   668 => x"fe01abb7",
   669 => x"48c187e1",
   670 => x"cef28ef0",
   671 => x"5b5e0e87",
   672 => x"710e5d5c",
   673 => x"c7029b4b",
   674 => x"4da3c887",
   675 => x"87c5056d",
   676 => x"fdc048ff",
   677 => x"4ca3d087",
   678 => x"ffc7496c",
   679 => x"87d80599",
   680 => x"87c9026c",
   681 => x"49731ec1",
   682 => x"c487f3f6",
   683 => x"e6e4c286",
   684 => x"f849731e",
   685 => x"86c487c2",
   686 => x"aa6d4a6c",
   687 => x"ff87c404",
   688 => x"c187cf48",
   689 => x"49727ca2",
   690 => x"c299ffc7",
   691 => x"9781e6e4",
   692 => x"f6f04869",
   693 => x"1e731e87",
   694 => x"029b4b71",
   695 => x"c287e4c0",
   696 => x"735bd3f1",
   697 => x"c28ac24a",
   698 => x"49bfe6ec",
   699 => x"fff0c292",
   700 => x"807248bf",
   701 => x"58d7f1c2",
   702 => x"30c44871",
   703 => x"58f6ecc2",
   704 => x"c287edc0",
   705 => x"c248cff1",
   706 => x"78bfc3f1",
   707 => x"48d3f1c2",
   708 => x"bfc7f1c2",
   709 => x"eeecc278",
   710 => x"87c902bf",
   711 => x"bfe6ecc2",
   712 => x"c731c449",
   713 => x"cbf1c287",
   714 => x"31c449bf",
   715 => x"59f6ecc2",
   716 => x"0e87dcef",
   717 => x"0e5c5b5e",
   718 => x"4bc04a71",
   719 => x"c0029a72",
   720 => x"a2da87e1",
   721 => x"4b699f49",
   722 => x"bfeeecc2",
   723 => x"d487cf02",
   724 => x"699f49a2",
   725 => x"ffc04c49",
   726 => x"34d09cff",
   727 => x"4cc087c2",
   728 => x"73b34974",
   729 => x"87edfd49",
   730 => x"0e87e2ee",
   731 => x"5d5c5b5e",
   732 => x"7186f40e",
   733 => x"727ec04a",
   734 => x"87d8029a",
   735 => x"48e2e4c2",
   736 => x"e4c278c0",
   737 => x"f1c248da",
   738 => x"c278bfd3",
   739 => x"c248dee4",
   740 => x"78bfcff1",
   741 => x"48c3edc2",
   742 => x"ecc250c0",
   743 => x"c249bff2",
   744 => x"4abfe2e4",
   745 => x"c403aa71",
   746 => x"497287ca",
   747 => x"c00599cf",
   748 => x"f5c087ea",
   749 => x"e4c248c7",
   750 => x"c278bfda",
   751 => x"c21ee6e4",
   752 => x"49bfdae4",
   753 => x"48dae4c2",
   754 => x"7178a1c1",
   755 => x"87fddeff",
   756 => x"f5c086c4",
   757 => x"e4c248c3",
   758 => x"87cc78e6",
   759 => x"bfc3f5c0",
   760 => x"80e0c048",
   761 => x"58c7f5c0",
   762 => x"bfe2e4c2",
   763 => x"c280c148",
   764 => x"2758e6e4",
   765 => x"00000d43",
   766 => x"4dbf97bf",
   767 => x"e3c2029d",
   768 => x"ade5c387",
   769 => x"87dcc202",
   770 => x"bfc3f5c0",
   771 => x"49a3cb4b",
   772 => x"accf4c11",
   773 => x"87d2c105",
   774 => x"99df4975",
   775 => x"91cd89c1",
   776 => x"81f6ecc2",
   777 => x"124aa3c1",
   778 => x"4aa3c351",
   779 => x"a3c55112",
   780 => x"c751124a",
   781 => x"51124aa3",
   782 => x"124aa3c9",
   783 => x"4aa3ce51",
   784 => x"a3d05112",
   785 => x"d251124a",
   786 => x"51124aa3",
   787 => x"124aa3d4",
   788 => x"4aa3d651",
   789 => x"a3d85112",
   790 => x"dc51124a",
   791 => x"51124aa3",
   792 => x"124aa3de",
   793 => x"c07ec151",
   794 => x"497487fa",
   795 => x"c00599c8",
   796 => x"497487eb",
   797 => x"d10599d0",
   798 => x"0266dc87",
   799 => x"7387cbc0",
   800 => x"0f66dc49",
   801 => x"c0029870",
   802 => x"056e87d3",
   803 => x"c287c6c0",
   804 => x"c048f6ec",
   805 => x"c3f5c050",
   806 => x"e1c248bf",
   807 => x"c3edc287",
   808 => x"7e50c048",
   809 => x"bff2ecc2",
   810 => x"e2e4c249",
   811 => x"aa714abf",
   812 => x"87f6fb04",
   813 => x"bfd3f1c2",
   814 => x"87c8c005",
   815 => x"bfeeecc2",
   816 => x"87f8c102",
   817 => x"bfdee4c2",
   818 => x"87c7e949",
   819 => x"e4c24970",
   820 => x"a6c459e2",
   821 => x"dee4c248",
   822 => x"ecc278bf",
   823 => x"c002bfee",
   824 => x"66c487d8",
   825 => x"ffffcf49",
   826 => x"a999f8ff",
   827 => x"87c5c002",
   828 => x"e1c04cc0",
   829 => x"c04cc187",
   830 => x"66c487dc",
   831 => x"f8ffcf49",
   832 => x"c002a999",
   833 => x"a6c887c8",
   834 => x"c078c048",
   835 => x"a6c887c5",
   836 => x"c878c148",
   837 => x"9c744c66",
   838 => x"87e0c005",
   839 => x"c24966c4",
   840 => x"e6ecc289",
   841 => x"c2914abf",
   842 => x"4abffff0",
   843 => x"48dae4c2",
   844 => x"c278a172",
   845 => x"c048e2e4",
   846 => x"87def978",
   847 => x"8ef448c0",
   848 => x"0087c8e7",
   849 => x"ff000000",
   850 => x"53ffffff",
   851 => x"5c00000d",
   852 => x"4600000d",
   853 => x"32335441",
   854 => x"00202020",
   855 => x"31544146",
   856 => x"20202036",
   857 => x"f1c21e00",
   858 => x"dd48bfd8",
   859 => x"87c905a8",
   860 => x"87cdc2c1",
   861 => x"c84a4970",
   862 => x"48d4ff87",
   863 => x"6878ffc3",
   864 => x"2648724a",
   865 => x"f1c21e4f",
   866 => x"dd48bfd8",
   867 => x"87c605a8",
   868 => x"87d9c1c1",
   869 => x"d4ff87d9",
   870 => x"78ffc348",
   871 => x"c048d0ff",
   872 => x"d4ff78e1",
   873 => x"c278d448",
   874 => x"ff48d7f1",
   875 => x"2650bfd4",
   876 => x"d0ff1e4f",
   877 => x"78e0c048",
   878 => x"fe1e4f26",
   879 => x"497087e7",
   880 => x"87c60299",
   881 => x"05a9fbc0",
   882 => x"487187f1",
   883 => x"5e0e4f26",
   884 => x"710e5c5b",
   885 => x"fe4cc04b",
   886 => x"497087cb",
   887 => x"f9c00299",
   888 => x"a9ecc087",
   889 => x"87f2c002",
   890 => x"02a9fbc0",
   891 => x"cc87ebc0",
   892 => x"03acb766",
   893 => x"66d087c7",
   894 => x"7187c202",
   895 => x"02997153",
   896 => x"84c187c2",
   897 => x"7087defd",
   898 => x"cd029949",
   899 => x"a9ecc087",
   900 => x"c087c702",
   901 => x"ff05a9fb",
   902 => x"66d087d5",
   903 => x"c087c302",
   904 => x"ecc07b97",
   905 => x"87c405a9",
   906 => x"87c54a74",
   907 => x"0ac04a74",
   908 => x"c248728a",
   909 => x"264d2687",
   910 => x"264b264c",
   911 => x"e4fc1e4f",
   912 => x"4a497087",
   913 => x"04aaf0c0",
   914 => x"f9c087c9",
   915 => x"87c301aa",
   916 => x"c18af0c0",
   917 => x"c904aac1",
   918 => x"aadac187",
   919 => x"c087c301",
   920 => x"48728af7",
   921 => x"5e0e4f26",
   922 => x"710e5c5b",
   923 => x"4cd4ff4a",
   924 => x"e9c04972",
   925 => x"9b4b7087",
   926 => x"c187c202",
   927 => x"48d0ff8b",
   928 => x"d5c178c5",
   929 => x"c649737c",
   930 => x"c3e7c131",
   931 => x"484abf97",
   932 => x"7c70b071",
   933 => x"c448d0ff",
   934 => x"fe487378",
   935 => x"5e0e87d9",
   936 => x"0e5d5c5b",
   937 => x"4b7186f8",
   938 => x"fec07ec0",
   939 => x"49bf97c4",
   940 => x"eec00599",
   941 => x"49a3c887",
   942 => x"c1496997",
   943 => x"dd05a9c1",
   944 => x"49a3c987",
   945 => x"c1496997",
   946 => x"d105a9d2",
   947 => x"49a3ca87",
   948 => x"c1496997",
   949 => x"c505a9c3",
   950 => x"c248df87",
   951 => x"48c087e1",
   952 => x"fa87dcc2",
   953 => x"4cc087df",
   954 => x"97c4fec0",
   955 => x"a9c049bf",
   956 => x"fb87cf04",
   957 => x"84c187c4",
   958 => x"97c4fec0",
   959 => x"06ac49bf",
   960 => x"fec087f1",
   961 => x"02bf97c4",
   962 => x"d8f987cf",
   963 => x"99497087",
   964 => x"c087c602",
   965 => x"f105a9ec",
   966 => x"f94cc087",
   967 => x"4d7087c7",
   968 => x"c887c2f9",
   969 => x"fcf858a6",
   970 => x"c14a7087",
   971 => x"49a3c884",
   972 => x"ad496997",
   973 => x"c087c702",
   974 => x"c005adff",
   975 => x"a3c987e7",
   976 => x"49699749",
   977 => x"02a966c4",
   978 => x"c04887c7",
   979 => x"d405a8ff",
   980 => x"49a3ca87",
   981 => x"aa496997",
   982 => x"c087c602",
   983 => x"c405aaff",
   984 => x"d07ec187",
   985 => x"adecc087",
   986 => x"c087c602",
   987 => x"c405adfb",
   988 => x"c14cc087",
   989 => x"fe026e7e",
   990 => x"f4f887e1",
   991 => x"f8487487",
   992 => x"87f1fa8e",
   993 => x"5b5e0e00",
   994 => x"f80e5d5c",
   995 => x"ff4d7186",
   996 => x"1e754bd4",
   997 => x"49dcf1c2",
   998 => x"87e9dfff",
   999 => x"987086c4",
  1000 => x"87fbc402",
  1001 => x"bfc5e7c1",
  1002 => x"fa49757e",
  1003 => x"a8de87f8",
  1004 => x"87ebc005",
  1005 => x"f6c04975",
  1006 => x"987087e5",
  1007 => x"c287db02",
  1008 => x"1ebfc0f6",
  1009 => x"c049e1c0",
  1010 => x"c487f4f3",
  1011 => x"c3e7c186",
  1012 => x"c250c048",
  1013 => x"fe49ccf6",
  1014 => x"48c187eb",
  1015 => x"ff87c2c4",
  1016 => x"78c548d0",
  1017 => x"c07bd6c1",
  1018 => x"49a2754a",
  1019 => x"82c17b11",
  1020 => x"04aab7cb",
  1021 => x"4acc87f3",
  1022 => x"c17bffc3",
  1023 => x"b7e0c082",
  1024 => x"87f404aa",
  1025 => x"c448d0ff",
  1026 => x"7bffc378",
  1027 => x"d3c178c5",
  1028 => x"c47bc17b",
  1029 => x"c0486e78",
  1030 => x"c206a8b7",
  1031 => x"f1c287f0",
  1032 => x"6e4cbfe4",
  1033 => x"70887448",
  1034 => x"029c747e",
  1035 => x"c287fdc1",
  1036 => x"c44de6e4",
  1037 => x"c0c848a6",
  1038 => x"b7c08c78",
  1039 => x"87c603ac",
  1040 => x"78a4c0c8",
  1041 => x"f1c24cc0",
  1042 => x"49bf97d7",
  1043 => x"d10299d0",
  1044 => x"c21ec087",
  1045 => x"e149dcf1",
  1046 => x"86c487de",
  1047 => x"c04a4970",
  1048 => x"e4c287ee",
  1049 => x"f1c21ee6",
  1050 => x"cbe149dc",
  1051 => x"7086c487",
  1052 => x"d0ff4a49",
  1053 => x"78c5c848",
  1054 => x"157bd4c1",
  1055 => x"4866c47b",
  1056 => x"a6c888c1",
  1057 => x"05987058",
  1058 => x"ff87f0ff",
  1059 => x"78c448d0",
  1060 => x"c5059a72",
  1061 => x"c148c087",
  1062 => x"1ec187c7",
  1063 => x"49dcf1c2",
  1064 => x"87fadeff",
  1065 => x"9c7486c4",
  1066 => x"87c3fe05",
  1067 => x"b7c0486e",
  1068 => x"87d106a8",
  1069 => x"48dcf1c2",
  1070 => x"80d078c0",
  1071 => x"80f478c0",
  1072 => x"bfe8f1c2",
  1073 => x"c0486e78",
  1074 => x"fd01a8b7",
  1075 => x"d0ff87d0",
  1076 => x"c178c548",
  1077 => x"7bc07bd3",
  1078 => x"48c178c4",
  1079 => x"c087c2c0",
  1080 => x"268ef848",
  1081 => x"264c264d",
  1082 => x"0e4f264b",
  1083 => x"5d5c5b5e",
  1084 => x"4b711e0e",
  1085 => x"ab4d4cc0",
  1086 => x"87e8c004",
  1087 => x"1edefac0",
  1088 => x"c4029d75",
  1089 => x"c24ac087",
  1090 => x"724ac187",
  1091 => x"87dbe949",
  1092 => x"7e7086c4",
  1093 => x"056e84c1",
  1094 => x"4c7387c2",
  1095 => x"ac7385c1",
  1096 => x"87d8ff06",
  1097 => x"fe26486e",
  1098 => x"711e87f9",
  1099 => x"0566c44a",
  1100 => x"497287c5",
  1101 => x"2687cef9",
  1102 => x"5b5e0e4f",
  1103 => x"1e0e5d5c",
  1104 => x"de494c71",
  1105 => x"c4f2c291",
  1106 => x"9785714d",
  1107 => x"dcc1026d",
  1108 => x"f0f1c287",
  1109 => x"82744abf",
  1110 => x"cefe4972",
  1111 => x"6e7e7087",
  1112 => x"87f2c002",
  1113 => x"4bf8f1c2",
  1114 => x"49cb4a6e",
  1115 => x"87f8fcfe",
  1116 => x"93cb4b74",
  1117 => x"83d7e7c1",
  1118 => x"c6c183c4",
  1119 => x"49747bf1",
  1120 => x"87fccac1",
  1121 => x"e7c17b75",
  1122 => x"49bf97c4",
  1123 => x"f8f1c21e",
  1124 => x"87d6fe49",
  1125 => x"497486c4",
  1126 => x"87e4cac1",
  1127 => x"ccc149c0",
  1128 => x"f1c287c3",
  1129 => x"78c048d8",
  1130 => x"d9dd49c1",
  1131 => x"f2fc2687",
  1132 => x"616f4c87",
  1133 => x"676e6964",
  1134 => x"002e2e2e",
  1135 => x"5c5b5e0e",
  1136 => x"4a4b710e",
  1137 => x"bff0f1c2",
  1138 => x"fc497282",
  1139 => x"4c7087dd",
  1140 => x"87c4029c",
  1141 => x"87dbe549",
  1142 => x"48f0f1c2",
  1143 => x"49c178c0",
  1144 => x"fb87e3dc",
  1145 => x"5e0e87ff",
  1146 => x"0e5d5c5b",
  1147 => x"e4c286f4",
  1148 => x"4cc04de6",
  1149 => x"c048a6c4",
  1150 => x"f0f1c278",
  1151 => x"a9c049bf",
  1152 => x"87c1c106",
  1153 => x"48e6e4c2",
  1154 => x"f8c00298",
  1155 => x"defac087",
  1156 => x"0266c81e",
  1157 => x"a6c487c7",
  1158 => x"c578c048",
  1159 => x"48a6c487",
  1160 => x"66c478c1",
  1161 => x"87c3e549",
  1162 => x"4d7086c4",
  1163 => x"66c484c1",
  1164 => x"c880c148",
  1165 => x"f1c258a6",
  1166 => x"ac49bff0",
  1167 => x"7587c603",
  1168 => x"c8ff059d",
  1169 => x"754cc087",
  1170 => x"e0c3029d",
  1171 => x"defac087",
  1172 => x"0266c81e",
  1173 => x"a6cc87c7",
  1174 => x"c578c048",
  1175 => x"48a6cc87",
  1176 => x"66cc78c1",
  1177 => x"87c3e449",
  1178 => x"7e7086c4",
  1179 => x"e9c2026e",
  1180 => x"cb496e87",
  1181 => x"49699781",
  1182 => x"c10299d0",
  1183 => x"c6c187d6",
  1184 => x"49744afc",
  1185 => x"e7c191cb",
  1186 => x"797281d7",
  1187 => x"ffc381c8",
  1188 => x"de497451",
  1189 => x"c4f2c291",
  1190 => x"c285714d",
  1191 => x"c17d97c1",
  1192 => x"e0c049a5",
  1193 => x"f6ecc251",
  1194 => x"d202bf97",
  1195 => x"c284c187",
  1196 => x"ecc24ba5",
  1197 => x"49db4af6",
  1198 => x"87ecf7fe",
  1199 => x"cd87dbc1",
  1200 => x"51c049a5",
  1201 => x"a5c284c1",
  1202 => x"cb4a6e4b",
  1203 => x"d7f7fe49",
  1204 => x"87c6c187",
  1205 => x"4af9c4c1",
  1206 => x"91cb4974",
  1207 => x"81d7e7c1",
  1208 => x"ecc27972",
  1209 => x"02bf97f6",
  1210 => x"497487d8",
  1211 => x"84c191de",
  1212 => x"4bc4f2c2",
  1213 => x"ecc28371",
  1214 => x"49dd4af6",
  1215 => x"87e8f6fe",
  1216 => x"4b7487d8",
  1217 => x"f2c293de",
  1218 => x"a3cb83c4",
  1219 => x"c151c049",
  1220 => x"4a6e7384",
  1221 => x"f6fe49cb",
  1222 => x"66c487ce",
  1223 => x"c880c148",
  1224 => x"acc758a6",
  1225 => x"87c5c003",
  1226 => x"e0fc056e",
  1227 => x"f4487487",
  1228 => x"87eff68e",
  1229 => x"711e731e",
  1230 => x"91cb494b",
  1231 => x"81d7e7c1",
  1232 => x"c14aa1c8",
  1233 => x"1248c3e7",
  1234 => x"4aa1c950",
  1235 => x"48c4fec0",
  1236 => x"81ca5012",
  1237 => x"48c4e7c1",
  1238 => x"e7c15011",
  1239 => x"49bf97c4",
  1240 => x"f749c01e",
  1241 => x"f1c287c4",
  1242 => x"78de48d8",
  1243 => x"d5d649c1",
  1244 => x"f2f52687",
  1245 => x"4a711e87",
  1246 => x"c191cb49",
  1247 => x"c881d7e7",
  1248 => x"c2481181",
  1249 => x"c258dcf1",
  1250 => x"c048f0f1",
  1251 => x"d549c178",
  1252 => x"4f2687f4",
  1253 => x"c149c01e",
  1254 => x"2687cac4",
  1255 => x"99711e4f",
  1256 => x"c187d202",
  1257 => x"c048ece8",
  1258 => x"c180f750",
  1259 => x"c140f5cd",
  1260 => x"ce78d0e7",
  1261 => x"e8e8c187",
  1262 => x"c9e7c148",
  1263 => x"c180fc78",
  1264 => x"2678d4ce",
  1265 => x"5b5e0e4f",
  1266 => x"4c710e5c",
  1267 => x"c192cb4a",
  1268 => x"c882d7e7",
  1269 => x"a2c949a2",
  1270 => x"4b6b974b",
  1271 => x"4969971e",
  1272 => x"1282ca1e",
  1273 => x"f6e4c049",
  1274 => x"d449c087",
  1275 => x"497487d8",
  1276 => x"87ccc1c1",
  1277 => x"ecf38ef8",
  1278 => x"1e731e87",
  1279 => x"ff494b71",
  1280 => x"497387c3",
  1281 => x"f387fefe",
  1282 => x"731e87dd",
  1283 => x"c64b711e",
  1284 => x"db024aa3",
  1285 => x"028ac187",
  1286 => x"028a87d6",
  1287 => x"8a87dac1",
  1288 => x"87fcc002",
  1289 => x"e1c0028a",
  1290 => x"cb028a87",
  1291 => x"87dbc187",
  1292 => x"c0fd49c7",
  1293 => x"87dec187",
  1294 => x"bff0f1c2",
  1295 => x"87cbc102",
  1296 => x"c288c148",
  1297 => x"c158f4f1",
  1298 => x"f1c287c1",
  1299 => x"c002bff4",
  1300 => x"f1c287f9",
  1301 => x"c148bff0",
  1302 => x"f4f1c280",
  1303 => x"87ebc058",
  1304 => x"bff0f1c2",
  1305 => x"c289c649",
  1306 => x"c059f4f1",
  1307 => x"da03a9b7",
  1308 => x"f0f1c287",
  1309 => x"d278c048",
  1310 => x"f4f1c287",
  1311 => x"87cb02bf",
  1312 => x"bff0f1c2",
  1313 => x"c280c648",
  1314 => x"c058f4f1",
  1315 => x"87f6d149",
  1316 => x"fec04973",
  1317 => x"cef187ea",
  1318 => x"1e731e87",
  1319 => x"f1c24b71",
  1320 => x"78dd48d8",
  1321 => x"ddd149c0",
  1322 => x"c0497387",
  1323 => x"f087d1fe",
  1324 => x"5e0e87f5",
  1325 => x"0e5d5c5b",
  1326 => x"d886ccff",
  1327 => x"a6c859a6",
  1328 => x"c478c048",
  1329 => x"66c8c180",
  1330 => x"c180c478",
  1331 => x"f4f1c278",
  1332 => x"c278c148",
  1333 => x"48bfd8f1",
  1334 => x"cb05a8de",
  1335 => x"87c6f487",
  1336 => x"a6cc4970",
  1337 => x"87d0cf59",
  1338 => x"e387dae2",
  1339 => x"f4e187cc",
  1340 => x"d44c7087",
  1341 => x"fcc10566",
  1342 => x"66c4c187",
  1343 => x"7080c448",
  1344 => x"48a6c47e",
  1345 => x"7278bf6e",
  1346 => x"ede3c11e",
  1347 => x"4966c848",
  1348 => x"204aa1c8",
  1349 => x"05aa7141",
  1350 => x"511087f9",
  1351 => x"c4c14a26",
  1352 => x"ccc14866",
  1353 => x"bf6e78f4",
  1354 => x"7481c749",
  1355 => x"66c4c151",
  1356 => x"c181c849",
  1357 => x"66c4c151",
  1358 => x"c081c949",
  1359 => x"66c4c151",
  1360 => x"c081ca49",
  1361 => x"acfbc051",
  1362 => x"c187cf02",
  1363 => x"c81ed81e",
  1364 => x"c849bf66",
  1365 => x"87f6e181",
  1366 => x"c8c186c8",
  1367 => x"a8c04866",
  1368 => x"c887c701",
  1369 => x"78c148a6",
  1370 => x"c8c187ce",
  1371 => x"88c14866",
  1372 => x"c358a6d0",
  1373 => x"87c2e187",
  1374 => x"c248a6d8",
  1375 => x"029c7478",
  1376 => x"c887f1cc",
  1377 => x"ccc14866",
  1378 => x"cc03a866",
  1379 => x"a6dc87e6",
  1380 => x"c478c048",
  1381 => x"ff78c080",
  1382 => x"7087cadf",
  1383 => x"4866d44c",
  1384 => x"c705a8dd",
  1385 => x"a6e0c087",
  1386 => x"7866d448",
  1387 => x"05acd0c1",
  1388 => x"ff87ebc0",
  1389 => x"ff87eede",
  1390 => x"7087eade",
  1391 => x"acecc04c",
  1392 => x"ff87c605",
  1393 => x"7087f3df",
  1394 => x"acd0c14c",
  1395 => x"d087c805",
  1396 => x"80c14866",
  1397 => x"c158a6d4",
  1398 => x"ff02acd0",
  1399 => x"e4c087d5",
  1400 => x"66d448a6",
  1401 => x"66e0c078",
  1402 => x"66e4c048",
  1403 => x"d5ca05a8",
  1404 => x"a6e8c087",
  1405 => x"ff78c048",
  1406 => x"78c080dc",
  1407 => x"fbc04d74",
  1408 => x"dbc9028d",
  1409 => x"028dc987",
  1410 => x"8dc287db",
  1411 => x"87f7c102",
  1412 => x"c4028dc9",
  1413 => x"8dc487d8",
  1414 => x"87c1c102",
  1415 => x"c4028dc1",
  1416 => x"f5c887cc",
  1417 => x"4966c887",
  1418 => x"c4c191cb",
  1419 => x"a1c48166",
  1420 => x"717e6a4a",
  1421 => x"f9e3c11e",
  1422 => x"4966c448",
  1423 => x"204aa1cc",
  1424 => x"05aa7141",
  1425 => x"1087f8ff",
  1426 => x"c1492651",
  1427 => x"ff79d9d2",
  1428 => x"7087d2dc",
  1429 => x"48a6c44c",
  1430 => x"c3c878c1",
  1431 => x"48a6dc87",
  1432 => x"ff78f0c0",
  1433 => x"7087fedb",
  1434 => x"acecc04c",
  1435 => x"87c4c002",
  1436 => x"5ca6e0c0",
  1437 => x"02acecc0",
  1438 => x"dbff87cd",
  1439 => x"4c7087e7",
  1440 => x"05acecc0",
  1441 => x"c087f3ff",
  1442 => x"c002acec",
  1443 => x"dbff87c4",
  1444 => x"1ec087d3",
  1445 => x"66d01eca",
  1446 => x"c191cb49",
  1447 => x"714866cc",
  1448 => x"58a6cc80",
  1449 => x"c44866c8",
  1450 => x"58a6d080",
  1451 => x"49bf66cc",
  1452 => x"87dadcff",
  1453 => x"1ede1ec1",
  1454 => x"49bf66d4",
  1455 => x"87cedcff",
  1456 => x"497086d0",
  1457 => x"c08909c0",
  1458 => x"c059a6f0",
  1459 => x"c04866ec",
  1460 => x"eec006a8",
  1461 => x"66ecc087",
  1462 => x"03a8dd48",
  1463 => x"c487e4c0",
  1464 => x"c049bf66",
  1465 => x"c08166ec",
  1466 => x"ecc051e0",
  1467 => x"81c14966",
  1468 => x"81bf66c4",
  1469 => x"c051c1c2",
  1470 => x"c24966ec",
  1471 => x"bf66c481",
  1472 => x"6e51c081",
  1473 => x"f4ccc148",
  1474 => x"c8496e78",
  1475 => x"5166d881",
  1476 => x"81c9496e",
  1477 => x"6e5166d0",
  1478 => x"dc81ca49",
  1479 => x"66d85166",
  1480 => x"dc80c148",
  1481 => x"ec4858a6",
  1482 => x"c478c180",
  1483 => x"dcff87f2",
  1484 => x"497087cb",
  1485 => x"59a6f0c0",
  1486 => x"87c1dcff",
  1487 => x"e0c04970",
  1488 => x"66dc59a6",
  1489 => x"a8ecc048",
  1490 => x"87cac005",
  1491 => x"c048a6dc",
  1492 => x"c07866ec",
  1493 => x"d8ff87c4",
  1494 => x"66c887cb",
  1495 => x"c191cb49",
  1496 => x"714866c4",
  1497 => x"6e7e7080",
  1498 => x"6e82c84a",
  1499 => x"c081ca49",
  1500 => x"dc5166ec",
  1501 => x"81c14966",
  1502 => x"8966ecc0",
  1503 => x"307148c1",
  1504 => x"89c14970",
  1505 => x"c27a9771",
  1506 => x"49bfe0f5",
  1507 => x"2966ecc0",
  1508 => x"484a6a97",
  1509 => x"f4c09871",
  1510 => x"496e58a6",
  1511 => x"48a681c4",
  1512 => x"e4c07869",
  1513 => x"e0c04866",
  1514 => x"c002a866",
  1515 => x"a6dc87c8",
  1516 => x"c078c048",
  1517 => x"a6dc87c5",
  1518 => x"dc78c148",
  1519 => x"e0c01e66",
  1520 => x"4966cc1e",
  1521 => x"87c6d8ff",
  1522 => x"4c7086c8",
  1523 => x"06acb7c0",
  1524 => x"c487dbc1",
  1525 => x"80744866",
  1526 => x"c058a6c8",
  1527 => x"897449e0",
  1528 => x"c14b66c4",
  1529 => x"714af6e3",
  1530 => x"87fce2fe",
  1531 => x"c24866c4",
  1532 => x"58a6c880",
  1533 => x"4866e8c0",
  1534 => x"ecc080c1",
  1535 => x"f0c058a6",
  1536 => x"81c14966",
  1537 => x"c002a970",
  1538 => x"4dc087c5",
  1539 => x"c187c2c0",
  1540 => x"c21e754d",
  1541 => x"e0c049a4",
  1542 => x"70887148",
  1543 => x"66cc1e49",
  1544 => x"e9d6ff49",
  1545 => x"c086c887",
  1546 => x"ff01a8b7",
  1547 => x"e8c087c6",
  1548 => x"d1c00266",
  1549 => x"c9496e87",
  1550 => x"66e8c081",
  1551 => x"c1486e51",
  1552 => x"c078c5cf",
  1553 => x"496e87cc",
  1554 => x"51c281c9",
  1555 => x"cfc1486e",
  1556 => x"a6c478f9",
  1557 => x"c078c148",
  1558 => x"d5ff87c6",
  1559 => x"4c7087dc",
  1560 => x"c00266c4",
  1561 => x"66c887f5",
  1562 => x"a866cc48",
  1563 => x"87cbc004",
  1564 => x"c14866c8",
  1565 => x"58a6cc80",
  1566 => x"cc87e0c0",
  1567 => x"88c14866",
  1568 => x"c058a6d0",
  1569 => x"c6c187d5",
  1570 => x"c8c005ac",
  1571 => x"4866d887",
  1572 => x"a6dc80c1",
  1573 => x"e1d4ff58",
  1574 => x"d04c7087",
  1575 => x"80c14866",
  1576 => x"7458a6d4",
  1577 => x"cbc0029c",
  1578 => x"4866c887",
  1579 => x"a866ccc1",
  1580 => x"87daf304",
  1581 => x"87f9d3ff",
  1582 => x"c74866c8",
  1583 => x"e5c003a8",
  1584 => x"f4f1c287",
  1585 => x"c878c048",
  1586 => x"91cb4966",
  1587 => x"8166c4c1",
  1588 => x"6a4aa1c4",
  1589 => x"7952c04a",
  1590 => x"c14866c8",
  1591 => x"58a6cc80",
  1592 => x"ff04a8c7",
  1593 => x"ccff87db",
  1594 => x"f6dfff8e",
  1595 => x"616f4c87",
  1596 => x"2e2a2064",
  1597 => x"203a0020",
  1598 => x"50494400",
  1599 => x"69775320",
  1600 => x"65686374",
  1601 => x"731e0073",
  1602 => x"9b4b711e",
  1603 => x"c287c602",
  1604 => x"c048f0f1",
  1605 => x"c21ec778",
  1606 => x"49bff0f1",
  1607 => x"d7e7c11e",
  1608 => x"d8f1c21e",
  1609 => x"c9ee49bf",
  1610 => x"c286cc87",
  1611 => x"49bfd8f1",
  1612 => x"7387eae9",
  1613 => x"87c8029b",
  1614 => x"49d7e7c1",
  1615 => x"87d2edc0",
  1616 => x"87e3deff",
  1617 => x"87c9c71e",
  1618 => x"f9fe49c1",
  1619 => x"e5e5fe87",
  1620 => x"02987087",
  1621 => x"ecfe87cd",
  1622 => x"987087fe",
  1623 => x"c187c402",
  1624 => x"c087c24a",
  1625 => x"059a724a",
  1626 => x"1ec087ce",
  1627 => x"49d5e6c1",
  1628 => x"87fcf8c0",
  1629 => x"87fe86c4",
  1630 => x"e6c11ec0",
  1631 => x"f8c049e0",
  1632 => x"1ec087ee",
  1633 => x"87c4fdc0",
  1634 => x"f8c04970",
  1635 => x"ffc287e2",
  1636 => x"268ef887",
  1637 => x"2044534f",
  1638 => x"6c696166",
  1639 => x"002e6465",
  1640 => x"746f6f42",
  1641 => x"2e676e69",
  1642 => x"1e002e2e",
  1643 => x"48f0f1c2",
  1644 => x"f1c278c0",
  1645 => x"78c048d8",
  1646 => x"c087c9fe",
  1647 => x"c087ecfc",
  1648 => x"004f2648",
  1649 => x"00000100",
  1650 => x"45208000",
  1651 => x"00746978",
  1652 => x"61422080",
  1653 => x"75006b63",
  1654 => x"84000013",
  1655 => x"0000002c",
  1656 => x"13750000",
  1657 => x"2ca20000",
  1658 => x"00000000",
  1659 => x"00137500",
  1660 => x"002cc000",
  1661 => x"00000000",
  1662 => x"00001375",
  1663 => x"00002cde",
  1664 => x"75000000",
  1665 => x"fc000013",
  1666 => x"0000002c",
  1667 => x"13750000",
  1668 => x"2d1a0000",
  1669 => x"00000000",
  1670 => x"00137500",
  1671 => x"002d3800",
  1672 => x"00000000",
  1673 => x"00001375",
  1674 => x"00000000",
  1675 => x"0a000000",
  1676 => x"00000014",
  1677 => x"00000000",
  1678 => x"fe1e0000",
  1679 => x"78c048f0",
  1680 => x"097909cd",
  1681 => x"1e1e4f26",
  1682 => x"7ebff0fe",
  1683 => x"4f262648",
  1684 => x"48f0fe1e",
  1685 => x"4f2678c1",
  1686 => x"48f0fe1e",
  1687 => x"4f2678c0",
  1688 => x"c04a711e",
  1689 => x"4f265252",
  1690 => x"5c5b5e0e",
  1691 => x"86f40e5d",
  1692 => x"6d974d71",
  1693 => x"4ca5c17e",
  1694 => x"c8486c97",
  1695 => x"486e58a6",
  1696 => x"05a866c4",
  1697 => x"48ff87c5",
  1698 => x"ff87e6c0",
  1699 => x"a5c287ca",
  1700 => x"4b6c9749",
  1701 => x"974ba371",
  1702 => x"6c974b6b",
  1703 => x"c1486e7e",
  1704 => x"58a6c880",
  1705 => x"a6cc98c7",
  1706 => x"7c977058",
  1707 => x"7387e1fe",
  1708 => x"268ef448",
  1709 => x"264c264d",
  1710 => x"0e4f264b",
  1711 => x"0e5c5b5e",
  1712 => x"4c7186f4",
  1713 => x"c34a66d8",
  1714 => x"a4c29aff",
  1715 => x"496c974b",
  1716 => x"7249a173",
  1717 => x"7e6c9751",
  1718 => x"80c1486e",
  1719 => x"c758a6c8",
  1720 => x"58a6cc98",
  1721 => x"8ef45470",
  1722 => x"1e87caff",
  1723 => x"87e8fd1e",
  1724 => x"494abfe0",
  1725 => x"99c0e0c0",
  1726 => x"7287cb02",
  1727 => x"d6f5c21e",
  1728 => x"87f7fe49",
  1729 => x"fdfc86c4",
  1730 => x"fd7e7087",
  1731 => x"262687c2",
  1732 => x"f5c21e4f",
  1733 => x"c7fd49d6",
  1734 => x"ebebc187",
  1735 => x"87dafc49",
  1736 => x"2687f7c3",
  1737 => x"5b5e0e4f",
  1738 => x"710e5d5c",
  1739 => x"d6f5c24d",
  1740 => x"87f4fc49",
  1741 => x"b7c04b70",
  1742 => x"c2c304ab",
  1743 => x"abf0c387",
  1744 => x"c187c905",
  1745 => x"c148c9f0",
  1746 => x"87e3c278",
  1747 => x"05abe0c3",
  1748 => x"f0c187c9",
  1749 => x"78c148cd",
  1750 => x"c187d4c2",
  1751 => x"02bfcdf0",
  1752 => x"c0c287c6",
  1753 => x"87c24ca3",
  1754 => x"f0c14c73",
  1755 => x"c002bfc9",
  1756 => x"497487e0",
  1757 => x"9129b7c4",
  1758 => x"81e9f1c1",
  1759 => x"9acf4a74",
  1760 => x"48c192c2",
  1761 => x"4a703072",
  1762 => x"4872baff",
  1763 => x"79709869",
  1764 => x"497487db",
  1765 => x"9129b7c4",
  1766 => x"81e9f1c1",
  1767 => x"9acf4a74",
  1768 => x"48c392c2",
  1769 => x"4a703072",
  1770 => x"70b06948",
  1771 => x"059d7579",
  1772 => x"ff87f0c0",
  1773 => x"e1c848d0",
  1774 => x"48d4ff78",
  1775 => x"f0c178c5",
  1776 => x"c302bfcd",
  1777 => x"78e0c387",
  1778 => x"bfc9f0c1",
  1779 => x"ff87c602",
  1780 => x"f0c348d4",
  1781 => x"48d4ff78",
  1782 => x"d0ff7873",
  1783 => x"78e1c848",
  1784 => x"c178e0c0",
  1785 => x"c048cdf0",
  1786 => x"c9f0c178",
  1787 => x"c278c048",
  1788 => x"f949d6f5",
  1789 => x"4b7087f2",
  1790 => x"03abb7c0",
  1791 => x"c087fefc",
  1792 => x"264d2648",
  1793 => x"264b264c",
  1794 => x"0000004f",
  1795 => x"00000000",
  1796 => x"4a711e00",
  1797 => x"87cdfc49",
  1798 => x"c01e4f26",
  1799 => x"c449724a",
  1800 => x"e9f1c191",
  1801 => x"c179c081",
  1802 => x"aab7d082",
  1803 => x"2687ee04",
  1804 => x"5b5e0e4f",
  1805 => x"710e5d5c",
  1806 => x"87dcf84d",
  1807 => x"b7c44a75",
  1808 => x"f1c1922a",
  1809 => x"4c7582e9",
  1810 => x"94c29ccf",
  1811 => x"744b496a",
  1812 => x"c29bc32b",
  1813 => x"70307448",
  1814 => x"74bcff4c",
  1815 => x"70987148",
  1816 => x"87ecf77a",
  1817 => x"d8fe4873",
  1818 => x"00000087",
  1819 => x"00000000",
  1820 => x"00000000",
  1821 => x"00000000",
  1822 => x"00000000",
  1823 => x"00000000",
  1824 => x"00000000",
  1825 => x"00000000",
  1826 => x"00000000",
  1827 => x"00000000",
  1828 => x"00000000",
  1829 => x"00000000",
  1830 => x"00000000",
  1831 => x"00000000",
  1832 => x"00000000",
  1833 => x"00000000",
  1834 => x"d0ff1e00",
  1835 => x"78e1c848",
  1836 => x"d4ff4871",
  1837 => x"66c47808",
  1838 => x"08d4ff48",
  1839 => x"1e4f2678",
  1840 => x"66c44a71",
  1841 => x"49721e49",
  1842 => x"ff87deff",
  1843 => x"e0c048d0",
  1844 => x"4f262678",
  1845 => x"711e731e",
  1846 => x"4966c84b",
  1847 => x"c14a731e",
  1848 => x"ff49a2e0",
  1849 => x"c42687d9",
  1850 => x"264d2687",
  1851 => x"264b264c",
  1852 => x"d4ff1e4f",
  1853 => x"7affc34a",
  1854 => x"c048d0ff",
  1855 => x"7ade78e1",
  1856 => x"bfe0f5c2",
  1857 => x"c848497a",
  1858 => x"717a7028",
  1859 => x"7028d048",
  1860 => x"d848717a",
  1861 => x"ff7a7028",
  1862 => x"e0c048d0",
  1863 => x"0e4f2678",
  1864 => x"5d5c5b5e",
  1865 => x"c24c710e",
  1866 => x"4dbfe0f5",
  1867 => x"71297449",
  1868 => x"9b66d04b",
  1869 => x"66d483c1",
  1870 => x"c204abb7",
  1871 => x"d04bc087",
  1872 => x"31744966",
  1873 => x"9975b9ff",
  1874 => x"32744a73",
  1875 => x"b0714872",
  1876 => x"58e4f5c2",
  1877 => x"2687dafe",
  1878 => x"264c264d",
  1879 => x"0e4f264b",
  1880 => x"5d5c5b5e",
  1881 => x"4c711e0e",
  1882 => x"4be4f5c2",
  1883 => x"f4c04ac0",
  1884 => x"c3cdfe49",
  1885 => x"c21e7487",
  1886 => x"fe49e4f5",
  1887 => x"c487c6e8",
  1888 => x"99497086",
  1889 => x"87eac002",
  1890 => x"4da61ec4",
  1891 => x"e4f5c21e",
  1892 => x"d4effe49",
  1893 => x"7086c887",
  1894 => x"87d60298",
  1895 => x"f7c14a75",
  1896 => x"4bc449e8",
  1897 => x"87c2cbfe",
  1898 => x"ca029870",
  1899 => x"c048c087",
  1900 => x"48c087ed",
  1901 => x"c087e8c0",
  1902 => x"c4c187f3",
  1903 => x"02987087",
  1904 => x"fcc087c8",
  1905 => x"05987087",
  1906 => x"f6c287f8",
  1907 => x"cc02bfc4",
  1908 => x"e0f5c287",
  1909 => x"c4f6c248",
  1910 => x"d4fc78bf",
  1911 => x"2648c187",
  1912 => x"4c264d26",
  1913 => x"4f264b26",
  1914 => x"4352415b",
  1915 => x"1ec01e00",
  1916 => x"49e4f5c2",
  1917 => x"87cfecfe",
  1918 => x"48fcf5c2",
  1919 => x"262678c0",
  1920 => x"5b5e0e4f",
  1921 => x"f40e5d5c",
  1922 => x"c27ec086",
  1923 => x"48bffcf5",
  1924 => x"03a8b7c3",
  1925 => x"f5c287d1",
  1926 => x"c148bffc",
  1927 => x"c0f6c280",
  1928 => x"48fbc058",
  1929 => x"c287d9c6",
  1930 => x"fe49e4f5",
  1931 => x"7087cef1",
  1932 => x"acb7c04c",
  1933 => x"4887c403",
  1934 => x"c287c5c6",
  1935 => x"4abffcf5",
  1936 => x"d8028ac3",
  1937 => x"028ac187",
  1938 => x"8a87c7c5",
  1939 => x"87f2c202",
  1940 => x"cfc1028a",
  1941 => x"c3028a87",
  1942 => x"d9c587de",
  1943 => x"c84dc087",
  1944 => x"4a755ca6",
  1945 => x"ffc192c4",
  1946 => x"f5c282de",
  1947 => x"84754cf8",
  1948 => x"494b6c97",
  1949 => x"97a3c14b",
  1950 => x"11816a7c",
  1951 => x"58a6cc48",
  1952 => x"c84866c4",
  1953 => x"c302a866",
  1954 => x"7c97c087",
  1955 => x"c70566c8",
  1956 => x"fcf5c287",
  1957 => x"78a5c448",
  1958 => x"b7c485c1",
  1959 => x"c1ff04ad",
  1960 => x"87d2c487",
  1961 => x"bfc8f6c2",
  1962 => x"a8b7c848",
  1963 => x"ca87cb01",
  1964 => x"87c602ac",
  1965 => x"c005accd",
  1966 => x"f6c287f3",
  1967 => x"c84bbfc8",
  1968 => x"d203abb7",
  1969 => x"ccf6c287",
  1970 => x"c0817349",
  1971 => x"83c151e0",
  1972 => x"04abb7c8",
  1973 => x"c287eeff",
  1974 => x"c148d4f6",
  1975 => x"cfc150d2",
  1976 => x"50cdc150",
  1977 => x"80e450c0",
  1978 => x"c9c378c3",
  1979 => x"c8f6c287",
  1980 => x"c14849bf",
  1981 => x"ccf6c280",
  1982 => x"a0c44858",
  1983 => x"c2517481",
  1984 => x"f0c087f4",
  1985 => x"da04acb7",
  1986 => x"b7f9c087",
  1987 => x"87d301ac",
  1988 => x"bfc0f6c2",
  1989 => x"7491ca49",
  1990 => x"8af0c04a",
  1991 => x"48c0f6c2",
  1992 => x"ca78a172",
  1993 => x"c6c002ac",
  1994 => x"05accd87",
  1995 => x"c287c7c2",
  1996 => x"c348fcf5",
  1997 => x"87fec178",
  1998 => x"acb7f0c0",
  1999 => x"c087db04",
  2000 => x"01acb7f9",
  2001 => x"c287d3c0",
  2002 => x"49bfc4f6",
  2003 => x"4a7491d0",
  2004 => x"c28af0c0",
  2005 => x"7248c4f6",
  2006 => x"c1c178a1",
  2007 => x"c004acb7",
  2008 => x"c6c187db",
  2009 => x"c001acb7",
  2010 => x"f6c287d3",
  2011 => x"d049bfc4",
  2012 => x"c04a7491",
  2013 => x"f6c28af7",
  2014 => x"a17248c4",
  2015 => x"02acca78",
  2016 => x"cd87c6c0",
  2017 => x"edc005ac",
  2018 => x"fcf5c287",
  2019 => x"c078c348",
  2020 => x"e2c087e4",
  2021 => x"c6c005ac",
  2022 => x"7efbc087",
  2023 => x"ca87d7c0",
  2024 => x"c6c002ac",
  2025 => x"05accd87",
  2026 => x"c287c9c0",
  2027 => x"c348fcf5",
  2028 => x"87c2c078",
  2029 => x"026e7e74",
  2030 => x"6e87d0f9",
  2031 => x"99ffc348",
  2032 => x"dbf88ef4",
  2033 => x"4e4f4387",
  2034 => x"4d003d46",
  2035 => x"4e00444f",
  2036 => x"00454d41",
  2037 => x"41464544",
  2038 => x"3d544c55",
  2039 => x"1fc50030",
  2040 => x"1fcb0000",
  2041 => x"1fcf0000",
  2042 => x"1fd40000",
  2043 => x"ff1e0000",
  2044 => x"c9c848d0",
  2045 => x"ff487178",
  2046 => x"267808d4",
  2047 => x"4a711e4f",
  2048 => x"ff87eb49",
  2049 => x"78c848d0",
  2050 => x"731e4f26",
  2051 => x"c24b711e",
  2052 => x"02bfe4f6",
  2053 => x"ebc287c3",
  2054 => x"48d0ff87",
  2055 => x"7378c9c8",
  2056 => x"b1e0c049",
  2057 => x"7148d4ff",
  2058 => x"d8f6c278",
  2059 => x"c878c048",
  2060 => x"87c50266",
  2061 => x"c249ffc3",
  2062 => x"c249c087",
  2063 => x"cc59e0f6",
  2064 => x"87c60266",
  2065 => x"4ad5d5c5",
  2066 => x"ffcf87c4",
  2067 => x"f6c24aff",
  2068 => x"f6c25ae4",
  2069 => x"78c148e4",
  2070 => x"4d2687c4",
  2071 => x"4b264c26",
  2072 => x"5e0e4f26",
  2073 => x"0e5d5c5b",
  2074 => x"f6c24a71",
  2075 => x"724cbfe0",
  2076 => x"87cb029a",
  2077 => x"c291c849",
  2078 => x"714bc0c0",
  2079 => x"c287c483",
  2080 => x"c04bc0c4",
  2081 => x"7449134d",
  2082 => x"dcf6c299",
  2083 => x"d4ffb9bf",
  2084 => x"c1787148",
  2085 => x"c8852cb7",
  2086 => x"e804adb7",
  2087 => x"d8f6c287",
  2088 => x"80c848bf",
  2089 => x"58dcf6c2",
  2090 => x"1e87effe",
  2091 => x"4b711e73",
  2092 => x"029a4a13",
  2093 => x"497287cb",
  2094 => x"1387e7fe",
  2095 => x"f5059a4a",
  2096 => x"87dafe87",
  2097 => x"d8f6c21e",
  2098 => x"f6c249bf",
  2099 => x"a1c148d8",
  2100 => x"b7c0c478",
  2101 => x"87db03a9",
  2102 => x"c248d4ff",
  2103 => x"78bfdcf6",
  2104 => x"bfd8f6c2",
  2105 => x"d8f6c249",
  2106 => x"78a1c148",
  2107 => x"a9b7c0c4",
  2108 => x"ff87e504",
  2109 => x"78c848d0",
  2110 => x"48e4f6c2",
  2111 => x"4f2678c0",
  2112 => x"00000000",
  2113 => x"00000000",
  2114 => x"5f000000",
  2115 => x"0000005f",
  2116 => x"00030300",
  2117 => x"00000303",
  2118 => x"147f7f14",
  2119 => x"00147f7f",
  2120 => x"6b2e2400",
  2121 => x"00123a6b",
  2122 => x"18366a4c",
  2123 => x"0032566c",
  2124 => x"594f7e30",
  2125 => x"40683a77",
  2126 => x"07040000",
  2127 => x"00000003",
  2128 => x"3e1c0000",
  2129 => x"00004163",
  2130 => x"63410000",
  2131 => x"00001c3e",
  2132 => x"1c3e2a08",
  2133 => x"082a3e1c",
  2134 => x"3e080800",
  2135 => x"0008083e",
  2136 => x"e0800000",
  2137 => x"00000060",
  2138 => x"08080800",
  2139 => x"00080808",
  2140 => x"60000000",
  2141 => x"00000060",
  2142 => x"18306040",
  2143 => x"0103060c",
  2144 => x"597f3e00",
  2145 => x"003e7f4d",
  2146 => x"7f060400",
  2147 => x"0000007f",
  2148 => x"71634200",
  2149 => x"00464f59",
  2150 => x"49632200",
  2151 => x"00367f49",
  2152 => x"13161c18",
  2153 => x"00107f7f",
  2154 => x"45672700",
  2155 => x"00397d45",
  2156 => x"4b7e3c00",
  2157 => x"00307949",
  2158 => x"71010100",
  2159 => x"00070f79",
  2160 => x"497f3600",
  2161 => x"00367f49",
  2162 => x"494f0600",
  2163 => x"001e3f69",
  2164 => x"66000000",
  2165 => x"00000066",
  2166 => x"e6800000",
  2167 => x"00000066",
  2168 => x"14080800",
  2169 => x"00222214",
  2170 => x"14141400",
  2171 => x"00141414",
  2172 => x"14222200",
  2173 => x"00080814",
  2174 => x"51030200",
  2175 => x"00060f59",
  2176 => x"5d417f3e",
  2177 => x"001e1f55",
  2178 => x"097f7e00",
  2179 => x"007e7f09",
  2180 => x"497f7f00",
  2181 => x"00367f49",
  2182 => x"633e1c00",
  2183 => x"00414141",
  2184 => x"417f7f00",
  2185 => x"001c3e63",
  2186 => x"497f7f00",
  2187 => x"00414149",
  2188 => x"097f7f00",
  2189 => x"00010109",
  2190 => x"417f3e00",
  2191 => x"007a7b49",
  2192 => x"087f7f00",
  2193 => x"007f7f08",
  2194 => x"7f410000",
  2195 => x"0000417f",
  2196 => x"40602000",
  2197 => x"003f7f40",
  2198 => x"1c087f7f",
  2199 => x"00416336",
  2200 => x"407f7f00",
  2201 => x"00404040",
  2202 => x"0c067f7f",
  2203 => x"007f7f06",
  2204 => x"0c067f7f",
  2205 => x"007f7f18",
  2206 => x"417f3e00",
  2207 => x"003e7f41",
  2208 => x"097f7f00",
  2209 => x"00060f09",
  2210 => x"61417f3e",
  2211 => x"00407e7f",
  2212 => x"097f7f00",
  2213 => x"00667f19",
  2214 => x"4d6f2600",
  2215 => x"00327b59",
  2216 => x"7f010100",
  2217 => x"0001017f",
  2218 => x"407f3f00",
  2219 => x"003f7f40",
  2220 => x"703f0f00",
  2221 => x"000f3f70",
  2222 => x"18307f7f",
  2223 => x"007f7f30",
  2224 => x"1c366341",
  2225 => x"4163361c",
  2226 => x"7c060301",
  2227 => x"0103067c",
  2228 => x"4d597161",
  2229 => x"00414347",
  2230 => x"7f7f0000",
  2231 => x"00004141",
  2232 => x"0c060301",
  2233 => x"40603018",
  2234 => x"41410000",
  2235 => x"00007f7f",
  2236 => x"03060c08",
  2237 => x"00080c06",
  2238 => x"80808080",
  2239 => x"00808080",
  2240 => x"03000000",
  2241 => x"00000407",
  2242 => x"54742000",
  2243 => x"00787c54",
  2244 => x"447f7f00",
  2245 => x"00387c44",
  2246 => x"447c3800",
  2247 => x"00004444",
  2248 => x"447c3800",
  2249 => x"007f7f44",
  2250 => x"547c3800",
  2251 => x"00185c54",
  2252 => x"7f7e0400",
  2253 => x"00000505",
  2254 => x"a4bc1800",
  2255 => x"007cfca4",
  2256 => x"047f7f00",
  2257 => x"00787c04",
  2258 => x"3d000000",
  2259 => x"0000407d",
  2260 => x"80808000",
  2261 => x"00007dfd",
  2262 => x"107f7f00",
  2263 => x"00446c38",
  2264 => x"3f000000",
  2265 => x"0000407f",
  2266 => x"180c7c7c",
  2267 => x"00787c0c",
  2268 => x"047c7c00",
  2269 => x"00787c04",
  2270 => x"447c3800",
  2271 => x"00387c44",
  2272 => x"24fcfc00",
  2273 => x"00183c24",
  2274 => x"243c1800",
  2275 => x"00fcfc24",
  2276 => x"047c7c00",
  2277 => x"00080c04",
  2278 => x"545c4800",
  2279 => x"00207454",
  2280 => x"7f3f0400",
  2281 => x"00004444",
  2282 => x"407c3c00",
  2283 => x"007c7c40",
  2284 => x"603c1c00",
  2285 => x"001c3c60",
  2286 => x"30607c3c",
  2287 => x"003c7c60",
  2288 => x"10386c44",
  2289 => x"00446c38",
  2290 => x"e0bc1c00",
  2291 => x"001c3c60",
  2292 => x"74644400",
  2293 => x"00444c5c",
  2294 => x"3e080800",
  2295 => x"00414177",
  2296 => x"7f000000",
  2297 => x"0000007f",
  2298 => x"77414100",
  2299 => x"0008083e",
  2300 => x"03010102",
  2301 => x"00010202",
  2302 => x"7f7f7f7f",
  2303 => x"007f7f7f",
  2304 => x"1c1c0808",
  2305 => x"7f7f3e3e",
  2306 => x"3e3e7f7f",
  2307 => x"08081c1c",
  2308 => x"7c181000",
  2309 => x"0010187c",
  2310 => x"7c301000",
  2311 => x"0010307c",
  2312 => x"60603010",
  2313 => x"00061e78",
  2314 => x"183c6642",
  2315 => x"0042663c",
  2316 => x"c26a3878",
  2317 => x"00386cc6",
  2318 => x"60000060",
  2319 => x"00600000",
  2320 => x"5c5b5e0e",
  2321 => x"711e0e5d",
  2322 => x"f5f6c24c",
  2323 => x"4bc04dbf",
  2324 => x"ab741ec0",
  2325 => x"c487c702",
  2326 => x"78c048a6",
  2327 => x"a6c487c5",
  2328 => x"c478c148",
  2329 => x"49731e66",
  2330 => x"c887dfee",
  2331 => x"49e0c086",
  2332 => x"c487efef",
  2333 => x"496a4aa5",
  2334 => x"f187f0f0",
  2335 => x"85cb87c6",
  2336 => x"b7c883c1",
  2337 => x"c7ff04ab",
  2338 => x"4d262687",
  2339 => x"4b264c26",
  2340 => x"711e4f26",
  2341 => x"f9f6c24a",
  2342 => x"f9f6c25a",
  2343 => x"4978c748",
  2344 => x"2687ddfe",
  2345 => x"1e731e4f",
  2346 => x"b7c04a71",
  2347 => x"87d303aa",
  2348 => x"bfc5e0c2",
  2349 => x"c187c405",
  2350 => x"c087c24b",
  2351 => x"c9e0c24b",
  2352 => x"c287c45b",
  2353 => x"c25ac9e0",
  2354 => x"4abfc5e0",
  2355 => x"c0c19ac1",
  2356 => x"e8ec49a2",
  2357 => x"c248fc87",
  2358 => x"78bfc5e0",
  2359 => x"1e87effe",
  2360 => x"66c44a71",
  2361 => x"ff49721e",
  2362 => x"2687e9df",
  2363 => x"c21e4f26",
  2364 => x"49bfc5e0",
  2365 => x"87d9dcff",
  2366 => x"48edf6c2",
  2367 => x"c278bfe8",
  2368 => x"ec48e9f6",
  2369 => x"f6c278bf",
  2370 => x"494abfed",
  2371 => x"c899ffc3",
  2372 => x"48722ab7",
  2373 => x"f6c2b071",
  2374 => x"4f2658f5",
  2375 => x"5c5b5e0e",
  2376 => x"4b710e5d",
  2377 => x"c287c7ff",
  2378 => x"c048e8f6",
  2379 => x"ff497350",
  2380 => x"7087fedb",
  2381 => x"9cc24c49",
  2382 => x"cb49eecb",
  2383 => x"497087cf",
  2384 => x"e8f6c24d",
  2385 => x"c105bf97",
  2386 => x"66d087e4",
  2387 => x"f1f6c249",
  2388 => x"d70599bf",
  2389 => x"4966d487",
  2390 => x"bfe9f6c2",
  2391 => x"87cc0599",
  2392 => x"dbff4973",
  2393 => x"987087cb",
  2394 => x"87c2c102",
  2395 => x"fdfd4cc1",
  2396 => x"ca497587",
  2397 => x"987087e3",
  2398 => x"c287c602",
  2399 => x"c148e8f6",
  2400 => x"e8f6c250",
  2401 => x"c005bf97",
  2402 => x"f6c287e4",
  2403 => x"d049bff1",
  2404 => x"ff059966",
  2405 => x"f6c287d6",
  2406 => x"d449bfe9",
  2407 => x"ff059966",
  2408 => x"497387ca",
  2409 => x"87c9daff",
  2410 => x"fe059870",
  2411 => x"487487fe",
  2412 => x"0e87d7fb",
  2413 => x"5d5c5b5e",
  2414 => x"c086f40e",
  2415 => x"bfec4c4d",
  2416 => x"48a6c47e",
  2417 => x"bff5f6c2",
  2418 => x"c01ec178",
  2419 => x"fd49c71e",
  2420 => x"86c887ca",
  2421 => x"ce029870",
  2422 => x"fb49ff87",
  2423 => x"dac187c7",
  2424 => x"ccd9ff49",
  2425 => x"c24dc187",
  2426 => x"bf97e8f6",
  2427 => x"c987c302",
  2428 => x"f6c287c0",
  2429 => x"c24bbfed",
  2430 => x"05bfc5e0",
  2431 => x"c387ebc0",
  2432 => x"d8ff49fd",
  2433 => x"fac387eb",
  2434 => x"e4d8ff49",
  2435 => x"c3497387",
  2436 => x"1e7199ff",
  2437 => x"c6fb49c0",
  2438 => x"c8497387",
  2439 => x"1e7129b7",
  2440 => x"fafa49c1",
  2441 => x"c686c887",
  2442 => x"f6c287c1",
  2443 => x"9b4bbff1",
  2444 => x"c287dd02",
  2445 => x"49bfc1e0",
  2446 => x"7087dec7",
  2447 => x"87c40598",
  2448 => x"87d24bc0",
  2449 => x"c749e0c2",
  2450 => x"e0c287c3",
  2451 => x"87c658c5",
  2452 => x"48c1e0c2",
  2453 => x"497378c0",
  2454 => x"ce0599c2",
  2455 => x"49ebc387",
  2456 => x"87cdd7ff",
  2457 => x"99c24970",
  2458 => x"fb87c202",
  2459 => x"c149734c",
  2460 => x"87ce0599",
  2461 => x"ff49f4c3",
  2462 => x"7087f6d6",
  2463 => x"0299c249",
  2464 => x"4cfa87c2",
  2465 => x"99c84973",
  2466 => x"c387ce05",
  2467 => x"d6ff49f5",
  2468 => x"497087df",
  2469 => x"d50299c2",
  2470 => x"f9f6c287",
  2471 => x"87ca02bf",
  2472 => x"c288c148",
  2473 => x"c058fdf6",
  2474 => x"4cff87c2",
  2475 => x"49734dc1",
  2476 => x"ce0599c4",
  2477 => x"49f2c387",
  2478 => x"87f5d5ff",
  2479 => x"99c24970",
  2480 => x"c287dc02",
  2481 => x"7ebff9f6",
  2482 => x"a8b7c748",
  2483 => x"87cbc003",
  2484 => x"80c1486e",
  2485 => x"58fdf6c2",
  2486 => x"fe87c2c0",
  2487 => x"c34dc14c",
  2488 => x"d5ff49fd",
  2489 => x"497087cb",
  2490 => x"c00299c2",
  2491 => x"f6c287d5",
  2492 => x"c002bff9",
  2493 => x"f6c287c9",
  2494 => x"78c048f9",
  2495 => x"fd87c2c0",
  2496 => x"c34dc14c",
  2497 => x"d4ff49fa",
  2498 => x"497087e7",
  2499 => x"c00299c2",
  2500 => x"f6c287d9",
  2501 => x"c748bff9",
  2502 => x"c003a8b7",
  2503 => x"f6c287c9",
  2504 => x"78c748f9",
  2505 => x"fc87c2c0",
  2506 => x"c04dc14c",
  2507 => x"c003acb7",
  2508 => x"66c487d1",
  2509 => x"82d8c14a",
  2510 => x"c6c0026a",
  2511 => x"744b6a87",
  2512 => x"c00f7349",
  2513 => x"1ef0c31e",
  2514 => x"f749dac1",
  2515 => x"86c887ce",
  2516 => x"c0029870",
  2517 => x"a6c887e2",
  2518 => x"f9f6c248",
  2519 => x"66c878bf",
  2520 => x"c491cb49",
  2521 => x"80714866",
  2522 => x"bf6e7e70",
  2523 => x"87c8c002",
  2524 => x"c84bbf6e",
  2525 => x"0f734966",
  2526 => x"c0029d75",
  2527 => x"f6c287c8",
  2528 => x"f249bff9",
  2529 => x"e0c287fa",
  2530 => x"c002bfc9",
  2531 => x"c24987dd",
  2532 => x"987087c7",
  2533 => x"87d3c002",
  2534 => x"bff9f6c2",
  2535 => x"87e0f249",
  2536 => x"c0f449c0",
  2537 => x"c9e0c287",
  2538 => x"f478c048",
  2539 => x"87daf38e",
  2540 => x"5c5b5e0e",
  2541 => x"711e0e5d",
  2542 => x"f5f6c24c",
  2543 => x"cdc149bf",
  2544 => x"d1c14da1",
  2545 => x"747e6981",
  2546 => x"87cf029c",
  2547 => x"744ba5c4",
  2548 => x"f5f6c27b",
  2549 => x"f9f249bf",
  2550 => x"747b6e87",
  2551 => x"87c4059c",
  2552 => x"87c24bc0",
  2553 => x"49734bc1",
  2554 => x"d487faf2",
  2555 => x"87c70266",
  2556 => x"7087da49",
  2557 => x"c087c24a",
  2558 => x"cde0c24a",
  2559 => x"c9f2265a",
  2560 => x"00000087",
  2561 => x"00000000",
  2562 => x"00000000",
  2563 => x"4a711e00",
  2564 => x"49bfc8ff",
  2565 => x"2648a172",
  2566 => x"c8ff1e4f",
  2567 => x"c0fe89bf",
  2568 => x"c0c0c0c0",
  2569 => x"87c401a9",
  2570 => x"87c24ac0",
  2571 => x"48724ac1",
  2572 => x"c21e4f26",
  2573 => x"49bfdbe1",
  2574 => x"e1c2b9c1",
  2575 => x"d4ff59df",
  2576 => x"78ffc348",
  2577 => x"c048d0ff",
  2578 => x"d4ff78e1",
  2579 => x"c478c148",
  2580 => x"ff787131",
  2581 => x"e0c048d0",
  2582 => x"004f2678",
  2583 => x"0e000000",
  2584 => x"5d5c5b5e",
  2585 => x"e9f6c20e",
  2586 => x"e3c24abf",
  2587 => x"4c49bfc8",
  2588 => x"4d71bc72",
  2589 => x"87e0c7ff",
  2590 => x"49744bc0",
  2591 => x"c00299d0",
  2592 => x"d0ff87e7",
  2593 => x"78e1c848",
  2594 => x"c548d4ff",
  2595 => x"d0497578",
  2596 => x"87c30299",
  2597 => x"c278f0c3",
  2598 => x"7349f6e3",
  2599 => x"ff481181",
  2600 => x"ff7808d4",
  2601 => x"e0c048d0",
  2602 => x"2d2cc178",
  2603 => x"04abc883",
  2604 => x"ff87c7ff",
  2605 => x"c287d9c6",
  2606 => x"c248c8e3",
  2607 => x"78bfe9f6",
  2608 => x"4c264d26",
  2609 => x"4f264b26",
  2610 => x"00000000",
  2611 => x"c3e7c11e",
  2612 => x"c250de48",
  2613 => x"fe49dfe3",
  2614 => x"c087eada",
  2615 => x"504f2648",
  2616 => x"4d4b4355",
  2617 => x"41317e41",
  2618 => x"1e004352",
  2619 => x"fd87c4f3",
  2620 => x"87f887ed",
  2621 => x"1e164f26",
  2622 => x"362e2526",
  2623 => x"362e3e3d",
  others => ( x"00000000")
);

-- Xilinx Vivado attributes
attribute ram_style: string;
attribute ram_style of ram: signal is "block";

signal q_local : std_logic_vector((NB_COL * COL_WIDTH)-1 downto 0);

signal wea : std_logic_vector(NB_COL - 1 downto 0);

begin

	output:
	for i in 0 to NB_COL - 1 generate
		q((i + 1) * COL_WIDTH - 1 downto i * COL_WIDTH) <= q_local((i+1) * COL_WIDTH - 1 downto i * COL_WIDTH);
	end generate;
    
    -- Generate write enable signals
    -- The Block ram generator doesn't like it when the compare is done in the if statement it self.
    wea <= bytesel when we = '1' else (others => '0');

    process(clk)
    begin
        if rising_edge(clk) then
            q_local <= ram(to_integer(unsigned(addr)));
            for i in 0 to NB_COL - 1 loop
                if (wea(NB_COL-i-1) = '1') then
                    ram(to_integer(unsigned(addr)))((i + 1) * COL_WIDTH - 1 downto i * COL_WIDTH) <= d((i + 1) * COL_WIDTH - 1 downto i * COL_WIDTH);
                end if;
            end loop;
        end if;
    end process;

end arch;
