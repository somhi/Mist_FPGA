library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity controller_rom2 is
generic	(
	ADDR_WIDTH : integer := 8; -- ROM's address width (words, not bytes)
	COL_WIDTH  : integer := 8;  -- Column width (8bit -> byte)
	NB_COL     : integer := 4  -- Number of columns in memory
	);
port (
	clk : in std_logic;
	reset_n : in std_logic := '1';
	addr : in std_logic_vector(ADDR_WIDTH-1 downto 0);
	q : out std_logic_vector(31 downto 0);
	-- Allow writes - defaults supplied to simplify projects that don't need to write.
	d : in std_logic_vector(31 downto 0) := X"00000000";
	we : in std_logic := '0';
	bytesel : in std_logic_vector(3 downto 0) := "1111"
);
end entity;

architecture arch of controller_rom2 is

-- type word_t is std_logic_vector(31 downto 0);
type ram_type is array (0 to 2 ** ADDR_WIDTH - 1) of std_logic_vector(NB_COL * COL_WIDTH - 1 downto 0);

signal ram : ram_type :=
(

     0 => x"b7c492cf",
     1 => x"aab7752a",
     2 => x"4a87c103",
     3 => x"06aab774",
     4 => x"724a87c1",
     5 => x"87d8fd7b",
     6 => x"d8cdc21e",
     7 => x"f5e449bf",
     8 => x"ede6c287",
     9 => x"78bfe848",
    10 => x"48e9e6c2",
    11 => x"c278bfec",
    12 => x"4abfede6",
    13 => x"99ffc349",
    14 => x"722ab7c8",
    15 => x"c2b07148",
    16 => x"2658f5e6",
    17 => x"5b5e0e4f",
    18 => x"710e5d5c",
    19 => x"87c8ff4b",
    20 => x"48e8e6c2",
    21 => x"497350c0",
    22 => x"7087dbe4",
    23 => x"9cc24c49",
    24 => x"cb49eecb",
    25 => x"497087fa",
    26 => x"e8e6c24d",
    27 => x"c105bf97",
    28 => x"66d087e2",
    29 => x"f1e6c249",
    30 => x"d60599bf",
    31 => x"4966d487",
    32 => x"bfe9e6c2",
    33 => x"87cb0599",
    34 => x"e9e34973",
    35 => x"02987087",
    36 => x"c187c1c1",
    37 => x"87c0fe4c",
    38 => x"cfcb4975",
    39 => x"02987087",
    40 => x"e6c287c6",
    41 => x"50c148e8",
    42 => x"97e8e6c2",
    43 => x"e3c005bf",
    44 => x"f1e6c287",
    45 => x"66d049bf",
    46 => x"d6ff0599",
    47 => x"e9e6c287",
    48 => x"66d449bf",
    49 => x"caff0599",
    50 => x"e2497387",
    51 => x"987087e8",
    52 => x"87fffe05",
    53 => x"d7fa4874",
    54 => x"5b5e0e87",
    55 => x"f40e5d5c",
    56 => x"4c4dc086",
    57 => x"c47ebfec",
    58 => x"e6c248a6",
    59 => x"c178bff5",
    60 => x"c71ec01e",
    61 => x"87cdfd49",
    62 => x"987086c8",
    63 => x"ff87cd02",
    64 => x"87c7fa49",
    65 => x"e149dac1",
    66 => x"4dc187ec",
    67 => x"97e8e6c2",
    68 => x"87c302bf",
    69 => x"c287eec9",
    70 => x"4bbfede6",
    71 => x"bfd8cdc2",
    72 => x"87d9c105",
    73 => x"c848a6c4",
    74 => x"c278c0c0",
    75 => x"6e7eddd4",
    76 => x"6e49bf97",
    77 => x"7080c148",
    78 => x"f9e0717e",
    79 => x"02987087",
    80 => x"66c487c3",
    81 => x"4866c4b3",
    82 => x"c828b7c1",
    83 => x"987058a6",
    84 => x"87dbff05",
    85 => x"e049fdc3",
    86 => x"fac387dc",
    87 => x"87d6e049",
    88 => x"ffc34973",
    89 => x"c01e7199",
    90 => x"87c6c949",
    91 => x"b7c84973",
    92 => x"c11e7129",
    93 => x"87fac849",
    94 => x"c1c686c8",
    95 => x"f1e6c287",
    96 => x"029b4bbf",
    97 => x"cdc287dd",
    98 => x"c749bfd4",
    99 => x"987087de",
   100 => x"c087c405",
   101 => x"c287d24b",
   102 => x"c3c749e0",
   103 => x"d8cdc287",
   104 => x"c287c658",
   105 => x"c048d4cd",
   106 => x"c2497378",
   107 => x"87ce0599",
   108 => x"ff49ebc3",
   109 => x"7087ffde",
   110 => x"0299c249",
   111 => x"4cfb87c2",
   112 => x"99c14973",
   113 => x"c387ce05",
   114 => x"deff49f4",
   115 => x"497087e8",
   116 => x"c20299c2",
   117 => x"734cfa87",
   118 => x"0599c849",
   119 => x"f5c387ce",
   120 => x"d1deff49",
   121 => x"c2497087",
   122 => x"87d50299",
   123 => x"bff9e6c2",
   124 => x"4887ca02",
   125 => x"e6c288c1",
   126 => x"c2c058fd",
   127 => x"c14cff87",
   128 => x"c449734d",
   129 => x"87ce0599",
   130 => x"ff49f2c3",
   131 => x"7087e7dd",
   132 => x"0299c249",
   133 => x"e6c287dc",
   134 => x"487ebff9",
   135 => x"03a8b7c7",
   136 => x"6e87cbc0",
   137 => x"c280c148",
   138 => x"c058fde6",
   139 => x"4cfe87c2",
   140 => x"fdc34dc1",
   141 => x"fddcff49",
   142 => x"c2497087",
   143 => x"d5c00299",
   144 => x"f9e6c287",
   145 => x"c9c002bf",
   146 => x"f9e6c287",
   147 => x"c078c048",
   148 => x"4cfd87c2",
   149 => x"fac34dc1",
   150 => x"d9dcff49",
   151 => x"c2497087",
   152 => x"d9c00299",
   153 => x"f9e6c287",
   154 => x"b7c748bf",
   155 => x"c9c003a8",
   156 => x"f9e6c287",
   157 => x"c078c748",
   158 => x"4cfc87c2",
   159 => x"b7c04dc1",
   160 => x"d1c003ac",
   161 => x"4a66c487",
   162 => x"6a82d8c1",
   163 => x"87c6c002",
   164 => x"49744b6a",
   165 => x"1ec00f73",
   166 => x"c11ef0c3",
   167 => x"e4f649da",
   168 => x"7086c887",
   169 => x"e2c00298",
   170 => x"48a6c887",
   171 => x"bff9e6c2",
   172 => x"4966c878",
   173 => x"66c491cb",
   174 => x"70807148",
   175 => x"02bf6e7e",
   176 => x"6e87c8c0",
   177 => x"66c84bbf",
   178 => x"750f7349",
   179 => x"c8c0029d",
   180 => x"f9e6c287",
   181 => x"cdf149bf",
   182 => x"dccdc287",
   183 => x"ddc002bf",
   184 => x"c7c24987",
   185 => x"02987087",
   186 => x"c287d3c0",
   187 => x"49bff9e6",
   188 => x"c087f3f0",
   189 => x"87d3f249",
   190 => x"48dccdc2",
   191 => x"8ef478c0",
   192 => x"0e87edf1",
   193 => x"5d5c5b5e",
   194 => x"4c711e0e",
   195 => x"bff5e6c2",
   196 => x"a1cdc149",
   197 => x"81d1c14d",
   198 => x"9c747e69",
   199 => x"c487cf02",
   200 => x"7b744ba5",
   201 => x"bff5e6c2",
   202 => x"87ccf149",
   203 => x"9c747b6e",
   204 => x"c087c405",
   205 => x"c187c24b",
   206 => x"f149734b",
   207 => x"66d487cd",
   208 => x"4987c702",
   209 => x"4a7087da",
   210 => x"4ac087c2",
   211 => x"5ae0cdc2",
   212 => x"87dcf026",
   213 => x"00000000",
   214 => x"00000000",
   215 => x"00000000",
   216 => x"ff4a711e",
   217 => x"7249bfc8",
   218 => x"4f2648a1",
   219 => x"bfc8ff1e",
   220 => x"c0c0fe89",
   221 => x"a9c0c0c0",
   222 => x"c087c401",
   223 => x"c187c24a",
   224 => x"2648724a",
   225 => x"cec21e4f",
   226 => x"c149bfee",
   227 => x"f2cec2b9",
   228 => x"48d4ff59",
   229 => x"ff78ffc3",
   230 => x"e1c048d0",
   231 => x"48d4ff78",
   232 => x"31c478c1",
   233 => x"d0ff7871",
   234 => x"78e0c048",
   235 => x"00004f26",
   236 => x"5e0e0000",
   237 => x"0e5d5c5b",
   238 => x"bfec4d71",
   239 => x"ff49c54b",
   240 => x"7087f3d6",
   241 => x"87c70598",
   242 => x"99c24973",
   243 => x"c287c702",
   244 => x"c248edd4",
   245 => x"49c678c0",
   246 => x"87dad6ff",
   247 => x"c7059870",
   248 => x"c4497387",
   249 => x"87c70299",
   250 => x"48edd4c2",
   251 => x"c478f0c0",
   252 => x"c1d6ff49",
   253 => x"05987087",
   254 => x"497387c7",
   255 => x"c60299c8",
   256 => x"edd4c287",
   257 => x"cc78cc48",
   258 => x"e9d5ff49",
   259 => x"05987087",
   260 => x"497387c7",
   261 => x"c60299d0",
   262 => x"edd4c287",
   263 => x"d078c848",
   264 => x"49751e66",
   265 => x"87f1d7ff",
   266 => x"bfedd4c2",
   267 => x"1e66d81e",
   268 => x"93c24b75",
   269 => x"94c84c75",
   270 => x"84fde6c2",
   271 => x"c4ee496c",
   272 => x"c27c7087",
   273 => x"1ebfedd4",
   274 => x"4966e0c0",
   275 => x"7129b7c2",
   276 => x"c293c41e",
   277 => x"6b83c1e7",
   278 => x"87e9ed49",
   279 => x"e6c27b70",
   280 => x"49751efd",
   281 => x"87ced7ff",
   282 => x"4d268ee8",
   283 => x"4b264c26",
   284 => x"731e4f26",
   285 => x"dfdcc11e",
   286 => x"c250c048",
   287 => x"c248f0d4",
   288 => x"c278c0c0",
   289 => x"48bfd4e6",
   290 => x"e6c2b0c1",
   291 => x"d7ff58d8",
   292 => x"d3c287d4",
   293 => x"e3fe49ee",
   294 => x"4b7087c2",
   295 => x"bfd4e6c2",
   296 => x"c298fe48",
   297 => x"ff58d8e6",
   298 => x"7387fbd6",
   299 => x"87c7059b",
   300 => x"48fad3c2",
   301 => x"c287f4c0",
   302 => x"48bfd4e6",
   303 => x"e6c2b0c1",
   304 => x"d6ff58d8",
   305 => x"d4c287e0",
   306 => x"78c148f0",
   307 => x"48dfdcc1",
   308 => x"d4c250c1",
   309 => x"e2fe49d1",
   310 => x"e6c287c2",
   311 => x"fe48bfd4",
   312 => x"d8e6c298",
   313 => x"fdd5ff58",
   314 => x"fe48c087",
   315 => x"455687c0",
   316 => x"45525443",
   317 => x"49422058",
   318 => x"4556004e",
   319 => x"45525443",
   320 => x"49422e58",
   321 => x"6f6e204e",
   322 => x"6f662074",
   323 => x"21646e75",
   324 => x"54554100",
   325 => x"4f4f424f",
   326 => x"43455654",
   327 => x"14125800",
   328 => x"1c1b1d11",
   329 => x"494a5923",
   330 => x"ebf2f541",
   331 => x"000080f4",
   332 => x"00008000",
  others => ( x"00000000")
);

-- Xilinx Vivado attributes
attribute ram_style: string;
attribute ram_style of ram: signal is "block";

signal q_local : std_logic_vector((NB_COL * COL_WIDTH)-1 downto 0);

signal wea : std_logic_vector(NB_COL - 1 downto 0);

begin

	output:
	for i in 0 to NB_COL - 1 generate
		q((i + 1) * COL_WIDTH - 1 downto i * COL_WIDTH) <= q_local((i+1) * COL_WIDTH - 1 downto i * COL_WIDTH);
	end generate;
    
    -- Generate write enable signals
    -- The Block ram generator doesn't like it when the compare is done in the if statement it self.
    wea <= bytesel when we = '1' else (others => '0');

    process(clk)
    begin
        if rising_edge(clk) then
            q_local <= ram(to_integer(unsigned(addr)));
            for i in 0 to NB_COL - 1 loop
                if (wea(NB_COL-i-1) = '1') then
                    ram(to_integer(unsigned(addr)))((i + 1) * COL_WIDTH - 1 downto i * COL_WIDTH) <= d((i + 1) * COL_WIDTH - 1 downto i * COL_WIDTH);
                end if;
            end loop;
        end if;
    end process;

end arch;
