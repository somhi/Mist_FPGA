library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity controller_rom2 is
generic	(
	ADDR_WIDTH : integer := 8; -- ROM's address width (words, not bytes)
	COL_WIDTH  : integer := 8;  -- Column width (8bit -> byte)
	NB_COL     : integer := 4  -- Number of columns in memory
	);
port (
	clk : in std_logic;
	reset_n : in std_logic := '1';
	addr : in std_logic_vector(ADDR_WIDTH-1 downto 0);
	q : out std_logic_vector(31 downto 0);
	-- Allow writes - defaults supplied to simplify projects that don't need to write.
	d : in std_logic_vector(31 downto 0) := X"00000000";
	we : in std_logic := '0';
	bytesel : in std_logic_vector(3 downto 0) := "1111"
);
end entity;

architecture arch of controller_rom2 is

-- type word_t is std_logic_vector(31 downto 0);
type ram_type is array (0 to 2 ** ADDR_WIDTH - 1) of std_logic_vector(NB_COL * COL_WIDTH - 1 downto 0);

signal ram : ram_type :=
(

     0 => x"4c554146",
     1 => x"00303d54",
     2 => x"00001fef",
     3 => x"00001ff5",
     4 => x"00001ff9",
     5 => x"00001ffe",
     6 => x"48d0ff1e",
     7 => x"7178c9c8",
     8 => x"08d4ff48",
     9 => x"1e4f2678",
    10 => x"eb494a71",
    11 => x"48d0ff87",
    12 => x"4f2678c8",
    13 => x"711e731e",
    14 => x"f0f9c24b",
    15 => x"87c302bf",
    16 => x"ff87ebc2",
    17 => x"c9c848d0",
    18 => x"c0497378",
    19 => x"d4ffb1e0",
    20 => x"c2787148",
    21 => x"c048e4f9",
    22 => x"0266c878",
    23 => x"ffc387c5",
    24 => x"c087c249",
    25 => x"ecf9c249",
    26 => x"0266cc59",
    27 => x"d5c587c6",
    28 => x"87c44ad5",
    29 => x"4affffcf",
    30 => x"5af0f9c2",
    31 => x"48f0f9c2",
    32 => x"87c478c1",
    33 => x"4c264d26",
    34 => x"4f264b26",
    35 => x"5c5b5e0e",
    36 => x"4a710e5d",
    37 => x"bfecf9c2",
    38 => x"029a724c",
    39 => x"c84987cb",
    40 => x"eac0c291",
    41 => x"c483714b",
    42 => x"eac4c287",
    43 => x"134dc04b",
    44 => x"c2997449",
    45 => x"b9bfe8f9",
    46 => x"7148d4ff",
    47 => x"2cb7c178",
    48 => x"adb7c885",
    49 => x"c287e804",
    50 => x"48bfe4f9",
    51 => x"f9c280c8",
    52 => x"effe58e8",
    53 => x"1e731e87",
    54 => x"4a134b71",
    55 => x"87cb029a",
    56 => x"e7fe4972",
    57 => x"9a4a1387",
    58 => x"fe87f505",
    59 => x"c21e87da",
    60 => x"49bfe4f9",
    61 => x"48e4f9c2",
    62 => x"c478a1c1",
    63 => x"03a9b7c0",
    64 => x"d4ff87db",
    65 => x"e8f9c248",
    66 => x"f9c278bf",
    67 => x"c249bfe4",
    68 => x"c148e4f9",
    69 => x"c0c478a1",
    70 => x"e504a9b7",
    71 => x"48d0ff87",
    72 => x"f9c278c8",
    73 => x"78c048f0",
    74 => x"00004f26",
    75 => x"00000000",
    76 => x"00000000",
    77 => x"005f5f00",
    78 => x"03000000",
    79 => x"03030003",
    80 => x"7f140000",
    81 => x"7f7f147f",
    82 => x"24000014",
    83 => x"3a6b6b2e",
    84 => x"6a4c0012",
    85 => x"566c1836",
    86 => x"7e300032",
    87 => x"3a77594f",
    88 => x"00004068",
    89 => x"00030704",
    90 => x"00000000",
    91 => x"41633e1c",
    92 => x"00000000",
    93 => x"1c3e6341",
    94 => x"2a080000",
    95 => x"3e1c1c3e",
    96 => x"0800082a",
    97 => x"083e3e08",
    98 => x"00000008",
    99 => x"0060e080",
   100 => x"08000000",
   101 => x"08080808",
   102 => x"00000008",
   103 => x"00606000",
   104 => x"60400000",
   105 => x"060c1830",
   106 => x"3e000103",
   107 => x"7f4d597f",
   108 => x"0400003e",
   109 => x"007f7f06",
   110 => x"42000000",
   111 => x"4f597163",
   112 => x"22000046",
   113 => x"7f494963",
   114 => x"1c180036",
   115 => x"7f7f1316",
   116 => x"27000010",
   117 => x"7d454567",
   118 => x"3c000039",
   119 => x"79494b7e",
   120 => x"01000030",
   121 => x"0f797101",
   122 => x"36000007",
   123 => x"7f49497f",
   124 => x"06000036",
   125 => x"3f69494f",
   126 => x"0000001e",
   127 => x"00666600",
   128 => x"00000000",
   129 => x"0066e680",
   130 => x"08000000",
   131 => x"22141408",
   132 => x"14000022",
   133 => x"14141414",
   134 => x"22000014",
   135 => x"08141422",
   136 => x"02000008",
   137 => x"0f595103",
   138 => x"7f3e0006",
   139 => x"1f555d41",
   140 => x"7e00001e",
   141 => x"7f09097f",
   142 => x"7f00007e",
   143 => x"7f49497f",
   144 => x"1c000036",
   145 => x"4141633e",
   146 => x"7f000041",
   147 => x"3e63417f",
   148 => x"7f00001c",
   149 => x"4149497f",
   150 => x"7f000041",
   151 => x"0109097f",
   152 => x"3e000001",
   153 => x"7b49417f",
   154 => x"7f00007a",
   155 => x"7f08087f",
   156 => x"0000007f",
   157 => x"417f7f41",
   158 => x"20000000",
   159 => x"7f404060",
   160 => x"7f7f003f",
   161 => x"63361c08",
   162 => x"7f000041",
   163 => x"4040407f",
   164 => x"7f7f0040",
   165 => x"7f060c06",
   166 => x"7f7f007f",
   167 => x"7f180c06",
   168 => x"3e00007f",
   169 => x"7f41417f",
   170 => x"7f00003e",
   171 => x"0f09097f",
   172 => x"7f3e0006",
   173 => x"7e7f6141",
   174 => x"7f000040",
   175 => x"7f19097f",
   176 => x"26000066",
   177 => x"7b594d6f",
   178 => x"01000032",
   179 => x"017f7f01",
   180 => x"3f000001",
   181 => x"7f40407f",
   182 => x"0f00003f",
   183 => x"3f70703f",
   184 => x"7f7f000f",
   185 => x"7f301830",
   186 => x"6341007f",
   187 => x"361c1c36",
   188 => x"03014163",
   189 => x"067c7c06",
   190 => x"71610103",
   191 => x"43474d59",
   192 => x"00000041",
   193 => x"41417f7f",
   194 => x"03010000",
   195 => x"30180c06",
   196 => x"00004060",
   197 => x"7f7f4141",
   198 => x"0c080000",
   199 => x"0c060306",
   200 => x"80800008",
   201 => x"80808080",
   202 => x"00000080",
   203 => x"04070300",
   204 => x"20000000",
   205 => x"7c545474",
   206 => x"7f000078",
   207 => x"7c44447f",
   208 => x"38000038",
   209 => x"4444447c",
   210 => x"38000000",
   211 => x"7f44447c",
   212 => x"3800007f",
   213 => x"5c54547c",
   214 => x"04000018",
   215 => x"05057f7e",
   216 => x"18000000",
   217 => x"fca4a4bc",
   218 => x"7f00007c",
   219 => x"7c04047f",
   220 => x"00000078",
   221 => x"407d3d00",
   222 => x"80000000",
   223 => x"7dfd8080",
   224 => x"7f000000",
   225 => x"6c38107f",
   226 => x"00000044",
   227 => x"407f3f00",
   228 => x"7c7c0000",
   229 => x"7c0c180c",
   230 => x"7c000078",
   231 => x"7c04047c",
   232 => x"38000078",
   233 => x"7c44447c",
   234 => x"fc000038",
   235 => x"3c2424fc",
   236 => x"18000018",
   237 => x"fc24243c",
   238 => x"7c0000fc",
   239 => x"0c04047c",
   240 => x"48000008",
   241 => x"7454545c",
   242 => x"04000020",
   243 => x"44447f3f",
   244 => x"3c000000",
   245 => x"7c40407c",
   246 => x"1c00007c",
   247 => x"3c60603c",
   248 => x"7c3c001c",
   249 => x"7c603060",
   250 => x"6c44003c",
   251 => x"6c381038",
   252 => x"1c000044",
   253 => x"3c60e0bc",
   254 => x"4400001c",
   255 => x"4c5c7464",
   256 => x"08000044",
   257 => x"41773e08",
   258 => x"00000041",
   259 => x"007f7f00",
   260 => x"41000000",
   261 => x"083e7741",
   262 => x"01020008",
   263 => x"02020301",
   264 => x"7f7f0001",
   265 => x"7f7f7f7f",
   266 => x"0808007f",
   267 => x"3e3e1c1c",
   268 => x"7f7f7f7f",
   269 => x"1c1c3e3e",
   270 => x"10000808",
   271 => x"187c7c18",
   272 => x"10000010",
   273 => x"307c7c30",
   274 => x"30100010",
   275 => x"1e786060",
   276 => x"66420006",
   277 => x"663c183c",
   278 => x"38780042",
   279 => x"6cc6c26a",
   280 => x"00600038",
   281 => x"00006000",
   282 => x"5e0e0060",
   283 => x"0e5d5c5b",
   284 => x"c24c711e",
   285 => x"4dbfc1fa",
   286 => x"1ec04bc0",
   287 => x"c702ab74",
   288 => x"48a6c487",
   289 => x"87c578c0",
   290 => x"c148a6c4",
   291 => x"1e66c478",
   292 => x"dfee4973",
   293 => x"c086c887",
   294 => x"efef49e0",
   295 => x"4aa5c487",
   296 => x"f0f0496a",
   297 => x"87c6f187",
   298 => x"83c185cb",
   299 => x"04abb7c8",
   300 => x"2687c7ff",
   301 => x"4c264d26",
   302 => x"4f264b26",
   303 => x"c24a711e",
   304 => x"c25ac5fa",
   305 => x"c748c5fa",
   306 => x"ddfe4978",
   307 => x"1e4f2687",
   308 => x"4a711e73",
   309 => x"03aab7c0",
   310 => x"e0c287d3",
   311 => x"c405bfef",
   312 => x"c24bc187",
   313 => x"c24bc087",
   314 => x"c45bf3e0",
   315 => x"f3e0c287",
   316 => x"efe0c25a",
   317 => x"9ac14abf",
   318 => x"49a2c0c1",
   319 => x"fc87e8ec",
   320 => x"efe0c248",
   321 => x"effe78bf",
   322 => x"4a711e87",
   323 => x"721e66c4",
   324 => x"dddfff49",
   325 => x"4f262687",
   326 => x"efe0c21e",
   327 => x"dcff49bf",
   328 => x"f9c287cd",
   329 => x"bfe848f9",
   330 => x"f5f9c278",
   331 => x"78bfec48",
   332 => x"bff9f9c2",
   333 => x"ffc3494a",
   334 => x"2ab7c899",
   335 => x"b0714872",
   336 => x"58c1fac2",
   337 => x"5e0e4f26",
   338 => x"0e5d5c5b",
   339 => x"c7ff4b71",
   340 => x"f4f9c287",
   341 => x"7350c048",
   342 => x"f2dbff49",
   343 => x"4c497087",
   344 => x"eecb9cc2",
   345 => x"87cfcb49",
   346 => x"c24d4970",
   347 => x"bf97f4f9",
   348 => x"87e4c105",
   349 => x"c24966d0",
   350 => x"99bffdf9",
   351 => x"d487d705",
   352 => x"f9c24966",
   353 => x"0599bff5",
   354 => x"497387cc",
   355 => x"87ffdaff",
   356 => x"c1029870",
   357 => x"4cc187c2",
   358 => x"7587fdfd",
   359 => x"87e3ca49",
   360 => x"c6029870",
   361 => x"f4f9c287",
   362 => x"c250c148",
   363 => x"bf97f4f9",
   364 => x"87e4c005",
   365 => x"bffdf9c2",
   366 => x"9966d049",
   367 => x"87d6ff05",
   368 => x"bff5f9c2",
   369 => x"9966d449",
   370 => x"87caff05",
   371 => x"d9ff4973",
   372 => x"987087fd",
   373 => x"87fefe05",
   374 => x"d7fb4874",
   375 => x"5b5e0e87",
   376 => x"f40e5d5c",
   377 => x"4c4dc086",
   378 => x"c47ebfec",
   379 => x"fac248a6",
   380 => x"c178bfc1",
   381 => x"c71ec01e",
   382 => x"87cafd49",
   383 => x"987086c8",
   384 => x"ff87ce02",
   385 => x"87c7fb49",
   386 => x"ff49dac1",
   387 => x"c187c0d9",
   388 => x"f4f9c24d",
   389 => x"c302bf97",
   390 => x"87c0c987",
   391 => x"bff9f9c2",
   392 => x"efe0c24b",
   393 => x"ebc005bf",
   394 => x"49fdc387",
   395 => x"87dfd8ff",
   396 => x"ff49fac3",
   397 => x"7387d8d8",
   398 => x"99ffc349",
   399 => x"49c01e71",
   400 => x"7387c6fb",
   401 => x"29b7c849",
   402 => x"49c11e71",
   403 => x"c887fafa",
   404 => x"87c1c686",
   405 => x"bffdf9c2",
   406 => x"dd029b4b",
   407 => x"ebe0c287",
   408 => x"dec749bf",
   409 => x"05987087",
   410 => x"4bc087c4",
   411 => x"e0c287d2",
   412 => x"87c3c749",
   413 => x"58efe0c2",
   414 => x"e0c287c6",
   415 => x"78c048eb",
   416 => x"99c24973",
   417 => x"c387ce05",
   418 => x"d7ff49eb",
   419 => x"497087c1",
   420 => x"c20299c2",
   421 => x"734cfb87",
   422 => x"0599c149",
   423 => x"f4c387ce",
   424 => x"ead6ff49",
   425 => x"c2497087",
   426 => x"87c20299",
   427 => x"49734cfa",
   428 => x"ce0599c8",
   429 => x"49f5c387",
   430 => x"87d3d6ff",
   431 => x"99c24970",
   432 => x"c287d502",
   433 => x"02bfc5fa",
   434 => x"c14887ca",
   435 => x"c9fac288",
   436 => x"87c2c058",
   437 => x"4dc14cff",
   438 => x"99c44973",
   439 => x"c387ce05",
   440 => x"d5ff49f2",
   441 => x"497087e9",
   442 => x"dc0299c2",
   443 => x"c5fac287",
   444 => x"c7487ebf",
   445 => x"c003a8b7",
   446 => x"486e87cb",
   447 => x"fac280c1",
   448 => x"c2c058c9",
   449 => x"c14cfe87",
   450 => x"49fdc34d",
   451 => x"87ffd4ff",
   452 => x"99c24970",
   453 => x"87d5c002",
   454 => x"bfc5fac2",
   455 => x"87c9c002",
   456 => x"48c5fac2",
   457 => x"c2c078c0",
   458 => x"c14cfd87",
   459 => x"49fac34d",
   460 => x"87dbd4ff",
   461 => x"99c24970",
   462 => x"87d9c002",
   463 => x"bfc5fac2",
   464 => x"a8b7c748",
   465 => x"87c9c003",
   466 => x"48c5fac2",
   467 => x"c2c078c7",
   468 => x"c14cfc87",
   469 => x"acb7c04d",
   470 => x"87d1c003",
   471 => x"c14a66c4",
   472 => x"026a82d8",
   473 => x"6a87c6c0",
   474 => x"7349744b",
   475 => x"c31ec00f",
   476 => x"dac11ef0",
   477 => x"87cef749",
   478 => x"987086c8",
   479 => x"87e2c002",
   480 => x"c248a6c8",
   481 => x"78bfc5fa",
   482 => x"cb4966c8",
   483 => x"4866c491",
   484 => x"7e708071",
   485 => x"c002bf6e",
   486 => x"bf6e87c8",
   487 => x"4966c84b",
   488 => x"9d750f73",
   489 => x"87c8c002",
   490 => x"bfc5fac2",
   491 => x"87faf249",
   492 => x"bff3e0c2",
   493 => x"87ddc002",
   494 => x"87c7c249",
   495 => x"c0029870",
   496 => x"fac287d3",
   497 => x"f249bfc5",
   498 => x"49c087e0",
   499 => x"c287c0f4",
   500 => x"c048f3e0",
   501 => x"f38ef478",
   502 => x"5e0e87da",
   503 => x"0e5d5c5b",
   504 => x"c24c711e",
   505 => x"49bfc1fa",
   506 => x"4da1cdc1",
   507 => x"6981d1c1",
   508 => x"029c747e",
   509 => x"a5c487cf",
   510 => x"c27b744b",
   511 => x"49bfc1fa",
   512 => x"6e87f9f2",
   513 => x"059c747b",
   514 => x"4bc087c4",
   515 => x"4bc187c2",
   516 => x"faf24973",
   517 => x"0266d487",
   518 => x"da4987c7",
   519 => x"c24a7087",
   520 => x"c24ac087",
   521 => x"265af7e0",
   522 => x"0087c9f2",
   523 => x"00000000",
   524 => x"00000000",
   525 => x"1e000000",
   526 => x"c8ff4a71",
   527 => x"a17249bf",
   528 => x"1e4f2648",
   529 => x"89bfc8ff",
   530 => x"c0c0c0fe",
   531 => x"01a9c0c0",
   532 => x"4ac087c4",
   533 => x"4ac187c2",
   534 => x"4f264872",
   535 => x"eae2c21e",
   536 => x"b9c149bf",
   537 => x"59eee2c2",
   538 => x"c348d4ff",
   539 => x"d0ff78ff",
   540 => x"78e1c048",
   541 => x"c148d4ff",
   542 => x"7131c478",
   543 => x"48d0ff78",
   544 => x"2678e0c0",
   545 => x"e2c21e4f",
   546 => x"f4c21ede",
   547 => x"fdfd49e8",
   548 => x"86c487df",
   549 => x"c3029870",
   550 => x"87c0ff87",
   551 => x"35314f26",
   552 => x"205a484b",
   553 => x"46432020",
   554 => x"00000047",
   555 => x"5e0e0000",
   556 => x"0e5d5c5b",
   557 => x"bff5f9c2",
   558 => x"d7e4c24a",
   559 => x"724c49bf",
   560 => x"ff4d71bc",
   561 => x"c087dec6",
   562 => x"d049744b",
   563 => x"e7c00299",
   564 => x"48d0ff87",
   565 => x"ff78e1c8",
   566 => x"78c548d4",
   567 => x"99d04975",
   568 => x"c387c302",
   569 => x"e7c278f0",
   570 => x"817349c4",
   571 => x"d4ff4811",
   572 => x"d0ff7808",
   573 => x"78e0c048",
   574 => x"832d2cc1",
   575 => x"ff04abc8",
   576 => x"c5ff87c7",
   577 => x"e4c287d7",
   578 => x"f9c248d7",
   579 => x"2678bff5",
   580 => x"264c264d",
   581 => x"004f264b",
   582 => x"1e000000",
   583 => x"4bc01e73",
   584 => x"48cce7c1",
   585 => x"1ec850de",
   586 => x"49c9fac2",
   587 => x"87ccd5fe",
   588 => x"1e7286c4",
   589 => x"48cde6c2",
   590 => x"49d1fac2",
   591 => x"204aa1c4",
   592 => x"05aa7141",
   593 => x"4a2687f9",
   594 => x"49d1e6c2",
   595 => x"87c2f9fd",
   596 => x"029a4a70",
   597 => x"fe4987c5",
   598 => x"7287ebc7",
   599 => x"dde6c21e",
   600 => x"d1fac248",
   601 => x"4aa1c449",
   602 => x"aa714120",
   603 => x"2687f905",
   604 => x"c9fac24a",
   605 => x"dcd9fe49",
   606 => x"05987087",
   607 => x"e6c287c4",
   608 => x"49c04be1",
   609 => x"87e0c5fe",
   610 => x"c6fe4873",
   611 => x"20202087",
   612 => x"544f4a00",
   613 => x"204f4745",
   614 => x"20202020",
   615 => x"43524100",
   616 => x"43524100",
   617 => x"746f6e20",
   618 => x"756f6620",
   619 => x"202e646e",
   620 => x"64616f4c",
   621 => x"43524120",
   622 => x"e0f01e00",
   623 => x"87eefb87",
   624 => x"4f2687f8",
   625 => x"25261e16",
   626 => x"3e3d362e",
  others => ( x"00000000")
);

-- Xilinx Vivado attributes
attribute ram_style: string;
attribute ram_style of ram: signal is "block";

signal q_local : std_logic_vector((NB_COL * COL_WIDTH)-1 downto 0);

signal wea : std_logic_vector(NB_COL - 1 downto 0);

begin

	output:
	for i in 0 to NB_COL - 1 generate
		q((i + 1) * COL_WIDTH - 1 downto i * COL_WIDTH) <= q_local((i+1) * COL_WIDTH - 1 downto i * COL_WIDTH);
	end generate;
    
    -- Generate write enable signals
    -- The Block ram generator doesn't like it when the compare is done in the if statement it self.
    wea <= bytesel when we = '1' else (others => '0');

    process(clk)
    begin
        if rising_edge(clk) then
            q_local <= ram(to_integer(unsigned(addr)));
            for i in 0 to NB_COL - 1 loop
                if (wea(NB_COL-i-1) = '1') then
                    ram(to_integer(unsigned(addr)))((i + 1) * COL_WIDTH - 1 downto i * COL_WIDTH) <= d((i + 1) * COL_WIDTH - 1 downto i * COL_WIDTH);
                end if;
            end loop;
        end if;
    end process;

end arch;
