
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity controller_rom is
generic
	(
		ADDR_WIDTH : integer := 15 -- Specify your actual ROM size to save LEs and unnecessary block RAM usage.
	);
port (
	clk : in std_logic;
	reset_n : in std_logic := '1';
	addr : in std_logic_vector(ADDR_WIDTH-1 downto 0);
	q : out std_logic_vector(31 downto 0);
	-- Allow writes - defaults supplied to simplify projects that don't need to write.
	d : in std_logic_vector(31 downto 0) := X"00000000";
	we : in std_logic := '0';
	bytesel : in std_logic_vector(3 downto 0) := "1111"
);
end entity;

architecture rtl of controller_rom is

	signal addr1 : integer range 0 to 2**ADDR_WIDTH-1;

	--  build up 2D array to hold the memory
	type word_t is array (0 to 3) of std_logic_vector(7 downto 0);
	type ram_t is array (0 to 2 ** ADDR_WIDTH - 1) of word_t;

	signal ram : ram_t:=
	(

     0 => (x"04",x"87",x"da",x"01"),
     1 => (x"58",x"0e",x"87",x"dd"),
     2 => (x"0e",x"5a",x"59",x"5e"),
     3 => (x"00",x"00",x"29",x"27"),
     4 => (x"4a",x"26",x"0f",x"00"),
     5 => (x"48",x"26",x"49",x"26"),
     6 => (x"08",x"26",x"80",x"ff"),
     7 => (x"00",x"2d",x"27",x"4f"),
     8 => (x"27",x"4f",x"00",x"00"),
     9 => (x"00",x"00",x"00",x"2a"),
    10 => (x"fd",x"00",x"4f",x"4f"),
    11 => (x"d0",x"e7",x"c2",x"87"),
    12 => (x"86",x"c0",x"c5",x"4e"),
    13 => (x"49",x"d0",x"e7",x"c2"),
    14 => (x"48",x"f4",x"d4",x"c2"),
    15 => (x"40",x"40",x"c0",x"89"),
    16 => (x"89",x"d0",x"40",x"40"),
    17 => (x"c1",x"87",x"f6",x"03"),
    18 => (x"00",x"87",x"fe",x"da"),
    19 => (x"1e",x"87",x"fc",x"98"),
    20 => (x"1e",x"73",x"1e",x"72"),
    21 => (x"02",x"11",x"48",x"12"),
    22 => (x"c3",x"4b",x"87",x"ca"),
    23 => (x"73",x"9b",x"98",x"df"),
    24 => (x"87",x"f0",x"02",x"88"),
    25 => (x"4a",x"26",x"4b",x"26"),
    26 => (x"73",x"1e",x"4f",x"26"),
    27 => (x"c1",x"1e",x"72",x"1e"),
    28 => (x"87",x"ca",x"04",x"8b"),
    29 => (x"02",x"11",x"48",x"12"),
    30 => (x"02",x"88",x"87",x"c4"),
    31 => (x"4a",x"26",x"87",x"f1"),
    32 => (x"4f",x"26",x"4b",x"26"),
    33 => (x"73",x"1e",x"74",x"1e"),
    34 => (x"c1",x"1e",x"72",x"1e"),
    35 => (x"87",x"d0",x"04",x"8b"),
    36 => (x"02",x"11",x"48",x"12"),
    37 => (x"c3",x"4c",x"87",x"ca"),
    38 => (x"74",x"9c",x"98",x"df"),
    39 => (x"87",x"eb",x"02",x"88"),
    40 => (x"4b",x"26",x"4a",x"26"),
    41 => (x"4f",x"26",x"4c",x"26"),
    42 => (x"81",x"48",x"73",x"1e"),
    43 => (x"c5",x"02",x"a9",x"73"),
    44 => (x"05",x"53",x"12",x"87"),
    45 => (x"4f",x"26",x"87",x"f6"),
    46 => (x"4a",x"66",x"c4",x"1e"),
    47 => (x"51",x"12",x"48",x"71"),
    48 => (x"26",x"87",x"fb",x"05"),
    49 => (x"4a",x"71",x"1e",x"4f"),
    50 => (x"48",x"49",x"66",x"c4"),
    51 => (x"a6",x"c8",x"88",x"c1"),
    52 => (x"02",x"99",x"71",x"58"),
    53 => (x"d4",x"ff",x"87",x"d6"),
    54 => (x"78",x"ff",x"c3",x"48"),
    55 => (x"66",x"c4",x"52",x"68"),
    56 => (x"88",x"c1",x"48",x"49"),
    57 => (x"71",x"58",x"a6",x"c8"),
    58 => (x"87",x"ea",x"05",x"99"),
    59 => (x"73",x"1e",x"4f",x"26"),
    60 => (x"4b",x"d4",x"ff",x"1e"),
    61 => (x"6b",x"7b",x"ff",x"c3"),
    62 => (x"7b",x"ff",x"c3",x"4a"),
    63 => (x"32",x"c8",x"49",x"6b"),
    64 => (x"ff",x"c3",x"b1",x"72"),
    65 => (x"c8",x"4a",x"6b",x"7b"),
    66 => (x"c3",x"b2",x"71",x"31"),
    67 => (x"49",x"6b",x"7b",x"ff"),
    68 => (x"b1",x"72",x"32",x"c8"),
    69 => (x"87",x"c4",x"48",x"71"),
    70 => (x"4c",x"26",x"4d",x"26"),
    71 => (x"4f",x"26",x"4b",x"26"),
    72 => (x"5c",x"5b",x"5e",x"0e"),
    73 => (x"4a",x"71",x"0e",x"5d"),
    74 => (x"72",x"4c",x"d4",x"ff"),
    75 => (x"99",x"ff",x"c3",x"49"),
    76 => (x"d4",x"c2",x"7c",x"71"),
    77 => (x"c8",x"05",x"bf",x"f4"),
    78 => (x"48",x"66",x"d0",x"87"),
    79 => (x"a6",x"d4",x"30",x"c9"),
    80 => (x"49",x"66",x"d0",x"58"),
    81 => (x"ff",x"c3",x"29",x"d8"),
    82 => (x"d0",x"7c",x"71",x"99"),
    83 => (x"29",x"d0",x"49",x"66"),
    84 => (x"71",x"99",x"ff",x"c3"),
    85 => (x"49",x"66",x"d0",x"7c"),
    86 => (x"ff",x"c3",x"29",x"c8"),
    87 => (x"d0",x"7c",x"71",x"99"),
    88 => (x"ff",x"c3",x"49",x"66"),
    89 => (x"72",x"7c",x"71",x"99"),
    90 => (x"c3",x"29",x"d0",x"49"),
    91 => (x"7c",x"71",x"99",x"ff"),
    92 => (x"f0",x"c9",x"4b",x"6c"),
    93 => (x"ff",x"c3",x"4d",x"ff"),
    94 => (x"87",x"d0",x"05",x"ab"),
    95 => (x"6c",x"7c",x"ff",x"c3"),
    96 => (x"02",x"8d",x"c1",x"4b"),
    97 => (x"ff",x"c3",x"87",x"c6"),
    98 => (x"87",x"f0",x"02",x"ab"),
    99 => (x"c7",x"fe",x"48",x"73"),
   100 => (x"49",x"c0",x"1e",x"87"),
   101 => (x"c3",x"48",x"d4",x"ff"),
   102 => (x"81",x"c1",x"78",x"ff"),
   103 => (x"a9",x"b7",x"c8",x"c3"),
   104 => (x"26",x"87",x"f1",x"04"),
   105 => (x"1e",x"73",x"1e",x"4f"),
   106 => (x"f8",x"c4",x"87",x"e7"),
   107 => (x"1e",x"c0",x"4b",x"df"),
   108 => (x"c1",x"f0",x"ff",x"c0"),
   109 => (x"e7",x"fd",x"49",x"f7"),
   110 => (x"c1",x"86",x"c4",x"87"),
   111 => (x"ea",x"c0",x"05",x"a8"),
   112 => (x"48",x"d4",x"ff",x"87"),
   113 => (x"c1",x"78",x"ff",x"c3"),
   114 => (x"c0",x"c0",x"c0",x"c0"),
   115 => (x"e1",x"c0",x"1e",x"c0"),
   116 => (x"49",x"e9",x"c1",x"f0"),
   117 => (x"c4",x"87",x"c9",x"fd"),
   118 => (x"05",x"98",x"70",x"86"),
   119 => (x"d4",x"ff",x"87",x"ca"),
   120 => (x"78",x"ff",x"c3",x"48"),
   121 => (x"87",x"cb",x"48",x"c1"),
   122 => (x"c1",x"87",x"e6",x"fe"),
   123 => (x"fd",x"fe",x"05",x"8b"),
   124 => (x"fc",x"48",x"c0",x"87"),
   125 => (x"73",x"1e",x"87",x"e6"),
   126 => (x"48",x"d4",x"ff",x"1e"),
   127 => (x"d3",x"78",x"ff",x"c3"),
   128 => (x"c0",x"1e",x"c0",x"4b"),
   129 => (x"c1",x"c1",x"f0",x"ff"),
   130 => (x"87",x"d4",x"fc",x"49"),
   131 => (x"98",x"70",x"86",x"c4"),
   132 => (x"ff",x"87",x"ca",x"05"),
   133 => (x"ff",x"c3",x"48",x"d4"),
   134 => (x"cb",x"48",x"c1",x"78"),
   135 => (x"87",x"f1",x"fd",x"87"),
   136 => (x"ff",x"05",x"8b",x"c1"),
   137 => (x"48",x"c0",x"87",x"db"),
   138 => (x"0e",x"87",x"f1",x"fb"),
   139 => (x"0e",x"5c",x"5b",x"5e"),
   140 => (x"fd",x"4c",x"d4",x"ff"),
   141 => (x"ea",x"c6",x"87",x"db"),
   142 => (x"f0",x"e1",x"c0",x"1e"),
   143 => (x"fb",x"49",x"c8",x"c1"),
   144 => (x"86",x"c4",x"87",x"de"),
   145 => (x"c8",x"02",x"a8",x"c1"),
   146 => (x"87",x"ea",x"fe",x"87"),
   147 => (x"e2",x"c1",x"48",x"c0"),
   148 => (x"87",x"da",x"fa",x"87"),
   149 => (x"ff",x"cf",x"49",x"70"),
   150 => (x"ea",x"c6",x"99",x"ff"),
   151 => (x"87",x"c8",x"02",x"a9"),
   152 => (x"c0",x"87",x"d3",x"fe"),
   153 => (x"87",x"cb",x"c1",x"48"),
   154 => (x"c0",x"7c",x"ff",x"c3"),
   155 => (x"f4",x"fc",x"4b",x"f1"),
   156 => (x"02",x"98",x"70",x"87"),
   157 => (x"c0",x"87",x"eb",x"c0"),
   158 => (x"f0",x"ff",x"c0",x"1e"),
   159 => (x"fa",x"49",x"fa",x"c1"),
   160 => (x"86",x"c4",x"87",x"de"),
   161 => (x"d9",x"05",x"98",x"70"),
   162 => (x"7c",x"ff",x"c3",x"87"),
   163 => (x"ff",x"c3",x"49",x"6c"),
   164 => (x"7c",x"7c",x"7c",x"7c"),
   165 => (x"02",x"99",x"c0",x"c1"),
   166 => (x"48",x"c1",x"87",x"c4"),
   167 => (x"48",x"c0",x"87",x"d5"),
   168 => (x"ab",x"c2",x"87",x"d1"),
   169 => (x"c0",x"87",x"c4",x"05"),
   170 => (x"c1",x"87",x"c8",x"48"),
   171 => (x"fd",x"fe",x"05",x"8b"),
   172 => (x"f9",x"48",x"c0",x"87"),
   173 => (x"73",x"1e",x"87",x"e4"),
   174 => (x"f4",x"d4",x"c2",x"1e"),
   175 => (x"c7",x"78",x"c1",x"48"),
   176 => (x"48",x"d0",x"ff",x"4b"),
   177 => (x"c8",x"fb",x"78",x"c2"),
   178 => (x"48",x"d0",x"ff",x"87"),
   179 => (x"1e",x"c0",x"78",x"c3"),
   180 => (x"c1",x"d0",x"e5",x"c0"),
   181 => (x"c7",x"f9",x"49",x"c0"),
   182 => (x"c1",x"86",x"c4",x"87"),
   183 => (x"87",x"c1",x"05",x"a8"),
   184 => (x"05",x"ab",x"c2",x"4b"),
   185 => (x"48",x"c0",x"87",x"c5"),
   186 => (x"c1",x"87",x"f9",x"c0"),
   187 => (x"d0",x"ff",x"05",x"8b"),
   188 => (x"87",x"f7",x"fc",x"87"),
   189 => (x"58",x"f8",x"d4",x"c2"),
   190 => (x"cd",x"05",x"98",x"70"),
   191 => (x"c0",x"1e",x"c1",x"87"),
   192 => (x"d0",x"c1",x"f0",x"ff"),
   193 => (x"87",x"d8",x"f8",x"49"),
   194 => (x"d4",x"ff",x"86",x"c4"),
   195 => (x"78",x"ff",x"c3",x"48"),
   196 => (x"c2",x"87",x"fc",x"c2"),
   197 => (x"ff",x"58",x"fc",x"d4"),
   198 => (x"78",x"c2",x"48",x"d0"),
   199 => (x"c3",x"48",x"d4",x"ff"),
   200 => (x"48",x"c1",x"78",x"ff"),
   201 => (x"0e",x"87",x"f5",x"f7"),
   202 => (x"5d",x"5c",x"5b",x"5e"),
   203 => (x"c0",x"4b",x"71",x"0e"),
   204 => (x"cd",x"ee",x"c5",x"4c"),
   205 => (x"d4",x"ff",x"4a",x"df"),
   206 => (x"78",x"ff",x"c3",x"48"),
   207 => (x"fe",x"c3",x"49",x"68"),
   208 => (x"fd",x"c0",x"05",x"a9"),
   209 => (x"73",x"4d",x"70",x"87"),
   210 => (x"87",x"cc",x"02",x"9b"),
   211 => (x"73",x"1e",x"66",x"d0"),
   212 => (x"87",x"f1",x"f5",x"49"),
   213 => (x"87",x"d6",x"86",x"c4"),
   214 => (x"c4",x"48",x"d0",x"ff"),
   215 => (x"ff",x"c3",x"78",x"d1"),
   216 => (x"48",x"66",x"d0",x"7d"),
   217 => (x"a6",x"d4",x"88",x"c1"),
   218 => (x"05",x"98",x"70",x"58"),
   219 => (x"d4",x"ff",x"87",x"f0"),
   220 => (x"78",x"ff",x"c3",x"48"),
   221 => (x"05",x"9b",x"73",x"78"),
   222 => (x"d0",x"ff",x"87",x"c5"),
   223 => (x"c1",x"78",x"d0",x"48"),
   224 => (x"8a",x"c1",x"4c",x"4a"),
   225 => (x"87",x"ee",x"fe",x"05"),
   226 => (x"cb",x"f6",x"48",x"74"),
   227 => (x"1e",x"73",x"1e",x"87"),
   228 => (x"4b",x"c0",x"4a",x"71"),
   229 => (x"c3",x"48",x"d4",x"ff"),
   230 => (x"d0",x"ff",x"78",x"ff"),
   231 => (x"78",x"c3",x"c4",x"48"),
   232 => (x"c3",x"48",x"d4",x"ff"),
   233 => (x"1e",x"72",x"78",x"ff"),
   234 => (x"c1",x"f0",x"ff",x"c0"),
   235 => (x"ef",x"f5",x"49",x"d1"),
   236 => (x"70",x"86",x"c4",x"87"),
   237 => (x"87",x"d2",x"05",x"98"),
   238 => (x"cc",x"1e",x"c0",x"c8"),
   239 => (x"e6",x"fd",x"49",x"66"),
   240 => (x"70",x"86",x"c4",x"87"),
   241 => (x"48",x"d0",x"ff",x"4b"),
   242 => (x"48",x"73",x"78",x"c2"),
   243 => (x"0e",x"87",x"cd",x"f5"),
   244 => (x"5d",x"5c",x"5b",x"5e"),
   245 => (x"c0",x"1e",x"c0",x"0e"),
   246 => (x"c9",x"c1",x"f0",x"ff"),
   247 => (x"87",x"c0",x"f5",x"49"),
   248 => (x"d4",x"c2",x"1e",x"d2"),
   249 => (x"fe",x"fc",x"49",x"fc"),
   250 => (x"c0",x"86",x"c8",x"87"),
   251 => (x"d2",x"84",x"c1",x"4c"),
   252 => (x"f8",x"04",x"ac",x"b7"),
   253 => (x"fc",x"d4",x"c2",x"87"),
   254 => (x"c3",x"49",x"bf",x"97"),
   255 => (x"c0",x"c1",x"99",x"c0"),
   256 => (x"e7",x"c0",x"05",x"a9"),
   257 => (x"c3",x"d5",x"c2",x"87"),
   258 => (x"d0",x"49",x"bf",x"97"),
   259 => (x"c4",x"d5",x"c2",x"31"),
   260 => (x"c8",x"4a",x"bf",x"97"),
   261 => (x"c2",x"b1",x"72",x"32"),
   262 => (x"bf",x"97",x"c5",x"d5"),
   263 => (x"4c",x"71",x"b1",x"4a"),
   264 => (x"ff",x"ff",x"ff",x"cf"),
   265 => (x"ca",x"84",x"c1",x"9c"),
   266 => (x"87",x"e7",x"c1",x"34"),
   267 => (x"97",x"c5",x"d5",x"c2"),
   268 => (x"31",x"c1",x"49",x"bf"),
   269 => (x"d5",x"c2",x"99",x"c6"),
   270 => (x"4a",x"bf",x"97",x"c6"),
   271 => (x"72",x"2a",x"b7",x"c7"),
   272 => (x"c1",x"d5",x"c2",x"b1"),
   273 => (x"4d",x"4a",x"bf",x"97"),
   274 => (x"d5",x"c2",x"9d",x"cf"),
   275 => (x"4a",x"bf",x"97",x"c2"),
   276 => (x"32",x"ca",x"9a",x"c3"),
   277 => (x"97",x"c3",x"d5",x"c2"),
   278 => (x"33",x"c2",x"4b",x"bf"),
   279 => (x"d5",x"c2",x"b2",x"73"),
   280 => (x"4b",x"bf",x"97",x"c4"),
   281 => (x"c6",x"9b",x"c0",x"c3"),
   282 => (x"b2",x"73",x"2b",x"b7"),
   283 => (x"48",x"c1",x"81",x"c2"),
   284 => (x"49",x"70",x"30",x"71"),
   285 => (x"30",x"75",x"48",x"c1"),
   286 => (x"4c",x"72",x"4d",x"70"),
   287 => (x"94",x"71",x"84",x"c1"),
   288 => (x"ad",x"b7",x"c0",x"c8"),
   289 => (x"c1",x"87",x"cc",x"06"),
   290 => (x"c8",x"2d",x"b7",x"34"),
   291 => (x"01",x"ad",x"b7",x"c0"),
   292 => (x"74",x"87",x"f4",x"ff"),
   293 => (x"87",x"c0",x"f2",x"48"),
   294 => (x"5c",x"5b",x"5e",x"0e"),
   295 => (x"86",x"f8",x"0e",x"5d"),
   296 => (x"48",x"e2",x"dd",x"c2"),
   297 => (x"d5",x"c2",x"78",x"c0"),
   298 => (x"49",x"c0",x"1e",x"da"),
   299 => (x"c4",x"87",x"de",x"fb"),
   300 => (x"05",x"98",x"70",x"86"),
   301 => (x"48",x"c0",x"87",x"c5"),
   302 => (x"c0",x"87",x"ce",x"c9"),
   303 => (x"c0",x"7e",x"c1",x"4d"),
   304 => (x"49",x"bf",x"c1",x"ee"),
   305 => (x"4a",x"d0",x"d6",x"c2"),
   306 => (x"ee",x"4b",x"c8",x"71"),
   307 => (x"98",x"70",x"87",x"dc"),
   308 => (x"c0",x"87",x"c2",x"05"),
   309 => (x"fd",x"ed",x"c0",x"7e"),
   310 => (x"d6",x"c2",x"49",x"bf"),
   311 => (x"c8",x"71",x"4a",x"ec"),
   312 => (x"87",x"c6",x"ee",x"4b"),
   313 => (x"c2",x"05",x"98",x"70"),
   314 => (x"6e",x"7e",x"c0",x"87"),
   315 => (x"87",x"fd",x"c0",x"02"),
   316 => (x"bf",x"e0",x"dc",x"c2"),
   317 => (x"d8",x"dd",x"c2",x"4d"),
   318 => (x"48",x"7e",x"bf",x"9f"),
   319 => (x"a8",x"ea",x"d6",x"c5"),
   320 => (x"c2",x"87",x"c7",x"05"),
   321 => (x"4d",x"bf",x"e0",x"dc"),
   322 => (x"48",x"6e",x"87",x"ce"),
   323 => (x"a8",x"d5",x"e9",x"ca"),
   324 => (x"c0",x"87",x"c5",x"02"),
   325 => (x"87",x"f1",x"c7",x"48"),
   326 => (x"1e",x"da",x"d5",x"c2"),
   327 => (x"ec",x"f9",x"49",x"75"),
   328 => (x"70",x"86",x"c4",x"87"),
   329 => (x"87",x"c5",x"05",x"98"),
   330 => (x"dc",x"c7",x"48",x"c0"),
   331 => (x"fd",x"ed",x"c0",x"87"),
   332 => (x"d6",x"c2",x"49",x"bf"),
   333 => (x"c8",x"71",x"4a",x"ec"),
   334 => (x"87",x"ee",x"ec",x"4b"),
   335 => (x"c8",x"05",x"98",x"70"),
   336 => (x"e2",x"dd",x"c2",x"87"),
   337 => (x"da",x"78",x"c1",x"48"),
   338 => (x"c1",x"ee",x"c0",x"87"),
   339 => (x"d6",x"c2",x"49",x"bf"),
   340 => (x"c8",x"71",x"4a",x"d0"),
   341 => (x"87",x"d2",x"ec",x"4b"),
   342 => (x"c0",x"02",x"98",x"70"),
   343 => (x"48",x"c0",x"87",x"c5"),
   344 => (x"c2",x"87",x"e6",x"c6"),
   345 => (x"bf",x"97",x"d8",x"dd"),
   346 => (x"a9",x"d5",x"c1",x"49"),
   347 => (x"87",x"cd",x"c0",x"05"),
   348 => (x"97",x"d9",x"dd",x"c2"),
   349 => (x"ea",x"c2",x"49",x"bf"),
   350 => (x"c5",x"c0",x"02",x"a9"),
   351 => (x"c6",x"48",x"c0",x"87"),
   352 => (x"d5",x"c2",x"87",x"c7"),
   353 => (x"7e",x"bf",x"97",x"da"),
   354 => (x"a8",x"e9",x"c3",x"48"),
   355 => (x"87",x"ce",x"c0",x"02"),
   356 => (x"eb",x"c3",x"48",x"6e"),
   357 => (x"c5",x"c0",x"02",x"a8"),
   358 => (x"c5",x"48",x"c0",x"87"),
   359 => (x"d5",x"c2",x"87",x"eb"),
   360 => (x"49",x"bf",x"97",x"e5"),
   361 => (x"cc",x"c0",x"05",x"99"),
   362 => (x"e6",x"d5",x"c2",x"87"),
   363 => (x"c2",x"49",x"bf",x"97"),
   364 => (x"c5",x"c0",x"02",x"a9"),
   365 => (x"c5",x"48",x"c0",x"87"),
   366 => (x"d5",x"c2",x"87",x"cf"),
   367 => (x"48",x"bf",x"97",x"e7"),
   368 => (x"58",x"de",x"dd",x"c2"),
   369 => (x"c1",x"48",x"4c",x"70"),
   370 => (x"e2",x"dd",x"c2",x"88"),
   371 => (x"e8",x"d5",x"c2",x"58"),
   372 => (x"75",x"49",x"bf",x"97"),
   373 => (x"e9",x"d5",x"c2",x"81"),
   374 => (x"c8",x"4a",x"bf",x"97"),
   375 => (x"7e",x"a1",x"72",x"32"),
   376 => (x"48",x"ef",x"e1",x"c2"),
   377 => (x"d5",x"c2",x"78",x"6e"),
   378 => (x"48",x"bf",x"97",x"ea"),
   379 => (x"c2",x"58",x"a6",x"c8"),
   380 => (x"02",x"bf",x"e2",x"dd"),
   381 => (x"c0",x"87",x"d4",x"c2"),
   382 => (x"49",x"bf",x"fd",x"ed"),
   383 => (x"4a",x"ec",x"d6",x"c2"),
   384 => (x"e9",x"4b",x"c8",x"71"),
   385 => (x"98",x"70",x"87",x"e4"),
   386 => (x"87",x"c5",x"c0",x"02"),
   387 => (x"f8",x"c3",x"48",x"c0"),
   388 => (x"da",x"dd",x"c2",x"87"),
   389 => (x"e2",x"c2",x"4c",x"bf"),
   390 => (x"d5",x"c2",x"5c",x"c3"),
   391 => (x"49",x"bf",x"97",x"ff"),
   392 => (x"d5",x"c2",x"31",x"c8"),
   393 => (x"4a",x"bf",x"97",x"fe"),
   394 => (x"d6",x"c2",x"49",x"a1"),
   395 => (x"4a",x"bf",x"97",x"c0"),
   396 => (x"a1",x"72",x"32",x"d0"),
   397 => (x"c1",x"d6",x"c2",x"49"),
   398 => (x"d8",x"4a",x"bf",x"97"),
   399 => (x"49",x"a1",x"72",x"32"),
   400 => (x"c2",x"91",x"66",x"c4"),
   401 => (x"81",x"bf",x"ef",x"e1"),
   402 => (x"59",x"f7",x"e1",x"c2"),
   403 => (x"97",x"c7",x"d6",x"c2"),
   404 => (x"32",x"c8",x"4a",x"bf"),
   405 => (x"97",x"c6",x"d6",x"c2"),
   406 => (x"4a",x"a2",x"4b",x"bf"),
   407 => (x"97",x"c8",x"d6",x"c2"),
   408 => (x"33",x"d0",x"4b",x"bf"),
   409 => (x"c2",x"4a",x"a2",x"73"),
   410 => (x"bf",x"97",x"c9",x"d6"),
   411 => (x"d8",x"9b",x"cf",x"4b"),
   412 => (x"4a",x"a2",x"73",x"33"),
   413 => (x"5a",x"fb",x"e1",x"c2"),
   414 => (x"bf",x"f7",x"e1",x"c2"),
   415 => (x"74",x"8a",x"c2",x"4a"),
   416 => (x"fb",x"e1",x"c2",x"92"),
   417 => (x"78",x"a1",x"72",x"48"),
   418 => (x"c2",x"87",x"ca",x"c1"),
   419 => (x"bf",x"97",x"ec",x"d5"),
   420 => (x"c2",x"31",x"c8",x"49"),
   421 => (x"bf",x"97",x"eb",x"d5"),
   422 => (x"c2",x"49",x"a1",x"4a"),
   423 => (x"c2",x"59",x"ea",x"dd"),
   424 => (x"49",x"bf",x"e6",x"dd"),
   425 => (x"ff",x"c7",x"31",x"c5"),
   426 => (x"c2",x"29",x"c9",x"81"),
   427 => (x"c2",x"59",x"c3",x"e2"),
   428 => (x"bf",x"97",x"f1",x"d5"),
   429 => (x"c2",x"32",x"c8",x"4a"),
   430 => (x"bf",x"97",x"f0",x"d5"),
   431 => (x"c4",x"4a",x"a2",x"4b"),
   432 => (x"82",x"6e",x"92",x"66"),
   433 => (x"5a",x"ff",x"e1",x"c2"),
   434 => (x"48",x"f7",x"e1",x"c2"),
   435 => (x"e1",x"c2",x"78",x"c0"),
   436 => (x"a1",x"72",x"48",x"f3"),
   437 => (x"c3",x"e2",x"c2",x"78"),
   438 => (x"f7",x"e1",x"c2",x"48"),
   439 => (x"e2",x"c2",x"78",x"bf"),
   440 => (x"e1",x"c2",x"48",x"c7"),
   441 => (x"c2",x"78",x"bf",x"fb"),
   442 => (x"02",x"bf",x"e2",x"dd"),
   443 => (x"74",x"87",x"c9",x"c0"),
   444 => (x"70",x"30",x"c4",x"48"),
   445 => (x"87",x"c9",x"c0",x"7e"),
   446 => (x"bf",x"ff",x"e1",x"c2"),
   447 => (x"70",x"30",x"c4",x"48"),
   448 => (x"e6",x"dd",x"c2",x"7e"),
   449 => (x"c1",x"78",x"6e",x"48"),
   450 => (x"26",x"8e",x"f8",x"48"),
   451 => (x"26",x"4c",x"26",x"4d"),
   452 => (x"0e",x"4f",x"26",x"4b"),
   453 => (x"5d",x"5c",x"5b",x"5e"),
   454 => (x"c2",x"4a",x"71",x"0e"),
   455 => (x"02",x"bf",x"e2",x"dd"),
   456 => (x"4b",x"72",x"87",x"cb"),
   457 => (x"4c",x"72",x"2b",x"c7"),
   458 => (x"c9",x"9c",x"ff",x"c1"),
   459 => (x"c8",x"4b",x"72",x"87"),
   460 => (x"c3",x"4c",x"72",x"2b"),
   461 => (x"e1",x"c2",x"9c",x"ff"),
   462 => (x"c0",x"83",x"bf",x"ef"),
   463 => (x"ab",x"bf",x"f9",x"ed"),
   464 => (x"c0",x"87",x"d9",x"02"),
   465 => (x"c2",x"5b",x"fd",x"ed"),
   466 => (x"73",x"1e",x"da",x"d5"),
   467 => (x"87",x"fd",x"f0",x"49"),
   468 => (x"98",x"70",x"86",x"c4"),
   469 => (x"c0",x"87",x"c5",x"05"),
   470 => (x"87",x"e6",x"c0",x"48"),
   471 => (x"bf",x"e2",x"dd",x"c2"),
   472 => (x"74",x"87",x"d2",x"02"),
   473 => (x"c2",x"91",x"c4",x"49"),
   474 => (x"69",x"81",x"da",x"d5"),
   475 => (x"ff",x"ff",x"cf",x"4d"),
   476 => (x"cb",x"9d",x"ff",x"ff"),
   477 => (x"c2",x"49",x"74",x"87"),
   478 => (x"da",x"d5",x"c2",x"91"),
   479 => (x"4d",x"69",x"9f",x"81"),
   480 => (x"c6",x"fe",x"48",x"75"),
   481 => (x"5b",x"5e",x"0e",x"87"),
   482 => (x"1e",x"0e",x"5d",x"5c"),
   483 => (x"1e",x"c0",x"4d",x"71"),
   484 => (x"c9",x"c8",x"49",x"c1"),
   485 => (x"70",x"86",x"c4",x"87"),
   486 => (x"c1",x"02",x"9c",x"4c"),
   487 => (x"dd",x"c2",x"87",x"c0"),
   488 => (x"49",x"75",x"4a",x"ea"),
   489 => (x"70",x"87",x"e8",x"e2"),
   490 => (x"f1",x"c0",x"02",x"98"),
   491 => (x"75",x"4a",x"74",x"87"),
   492 => (x"e3",x"4b",x"cb",x"49"),
   493 => (x"98",x"70",x"87",x"ce"),
   494 => (x"87",x"e2",x"c0",x"02"),
   495 => (x"9c",x"74",x"1e",x"c0"),
   496 => (x"c4",x"87",x"c7",x"02"),
   497 => (x"78",x"c0",x"48",x"a6"),
   498 => (x"a6",x"c4",x"87",x"c5"),
   499 => (x"c4",x"78",x"c1",x"48"),
   500 => (x"c9",x"c7",x"49",x"66"),
   501 => (x"70",x"86",x"c4",x"87"),
   502 => (x"ff",x"05",x"9c",x"4c"),
   503 => (x"48",x"74",x"87",x"c0"),
   504 => (x"87",x"e7",x"fc",x"26"),
   505 => (x"5c",x"5b",x"5e",x"0e"),
   506 => (x"71",x"1e",x"0e",x"5d"),
   507 => (x"c5",x"05",x"9b",x"4b"),
   508 => (x"c1",x"48",x"c0",x"87"),
   509 => (x"a3",x"c8",x"87",x"e5"),
   510 => (x"d4",x"7d",x"c0",x"4d"),
   511 => (x"87",x"c7",x"02",x"66"),
   512 => (x"bf",x"97",x"66",x"d4"),
   513 => (x"c0",x"87",x"c5",x"05"),
   514 => (x"87",x"cf",x"c1",x"48"),
   515 => (x"fd",x"49",x"66",x"d4"),
   516 => (x"4c",x"70",x"87",x"f3"),
   517 => (x"c0",x"c1",x"02",x"9c"),
   518 => (x"49",x"a4",x"dc",x"87"),
   519 => (x"a4",x"da",x"7d",x"69"),
   520 => (x"4a",x"a3",x"c4",x"49"),
   521 => (x"c2",x"7a",x"69",x"9f"),
   522 => (x"02",x"bf",x"e2",x"dd"),
   523 => (x"a4",x"d4",x"87",x"d2"),
   524 => (x"49",x"69",x"9f",x"49"),
   525 => (x"99",x"ff",x"ff",x"c0"),
   526 => (x"30",x"d0",x"48",x"71"),
   527 => (x"87",x"c2",x"7e",x"70"),
   528 => (x"49",x"6e",x"7e",x"c0"),
   529 => (x"70",x"80",x"6a",x"48"),
   530 => (x"cc",x"7b",x"c0",x"7a"),
   531 => (x"79",x"6a",x"49",x"a3"),
   532 => (x"c0",x"49",x"a3",x"d0"),
   533 => (x"c2",x"48",x"c1",x"79"),
   534 => (x"26",x"48",x"c0",x"87"),
   535 => (x"0e",x"87",x"ec",x"fa"),
   536 => (x"5d",x"5c",x"5b",x"5e"),
   537 => (x"9c",x"4c",x"71",x"0e"),
   538 => (x"87",x"ca",x"c1",x"02"),
   539 => (x"69",x"49",x"a4",x"c8"),
   540 => (x"87",x"c2",x"c1",x"02"),
   541 => (x"6c",x"4a",x"66",x"d0"),
   542 => (x"a6",x"d4",x"82",x"49"),
   543 => (x"4d",x"66",x"d0",x"5a"),
   544 => (x"de",x"dd",x"c2",x"b9"),
   545 => (x"ba",x"ff",x"4a",x"bf"),
   546 => (x"99",x"71",x"99",x"72"),
   547 => (x"87",x"e4",x"c0",x"02"),
   548 => (x"6b",x"4b",x"a4",x"c4"),
   549 => (x"87",x"fb",x"f9",x"49"),
   550 => (x"dd",x"c2",x"7b",x"70"),
   551 => (x"6c",x"49",x"bf",x"da"),
   552 => (x"75",x"7c",x"71",x"81"),
   553 => (x"de",x"dd",x"c2",x"b9"),
   554 => (x"ba",x"ff",x"4a",x"bf"),
   555 => (x"99",x"71",x"99",x"72"),
   556 => (x"87",x"dc",x"ff",x"05"),
   557 => (x"d2",x"f9",x"7c",x"75"),
   558 => (x"1e",x"73",x"1e",x"87"),
   559 => (x"02",x"9b",x"4b",x"71"),
   560 => (x"a3",x"c8",x"87",x"c7"),
   561 => (x"c5",x"05",x"69",x"49"),
   562 => (x"c0",x"48",x"c0",x"87"),
   563 => (x"e1",x"c2",x"87",x"f7"),
   564 => (x"c4",x"4a",x"bf",x"f3"),
   565 => (x"49",x"69",x"49",x"a3"),
   566 => (x"dd",x"c2",x"89",x"c2"),
   567 => (x"71",x"91",x"bf",x"da"),
   568 => (x"dd",x"c2",x"4a",x"a2"),
   569 => (x"6b",x"49",x"bf",x"de"),
   570 => (x"4a",x"a2",x"71",x"99"),
   571 => (x"5a",x"fd",x"ed",x"c0"),
   572 => (x"72",x"1e",x"66",x"c8"),
   573 => (x"87",x"d5",x"ea",x"49"),
   574 => (x"98",x"70",x"86",x"c4"),
   575 => (x"c0",x"87",x"c4",x"05"),
   576 => (x"c1",x"87",x"c2",x"48"),
   577 => (x"87",x"c7",x"f8",x"48"),
   578 => (x"71",x"1e",x"73",x"1e"),
   579 => (x"c0",x"02",x"9b",x"4b"),
   580 => (x"e2",x"c2",x"87",x"e4"),
   581 => (x"4a",x"73",x"5b",x"c7"),
   582 => (x"dd",x"c2",x"8a",x"c2"),
   583 => (x"92",x"49",x"bf",x"da"),
   584 => (x"bf",x"f3",x"e1",x"c2"),
   585 => (x"c2",x"80",x"72",x"48"),
   586 => (x"71",x"58",x"cb",x"e2"),
   587 => (x"c2",x"30",x"c4",x"48"),
   588 => (x"c0",x"58",x"ea",x"dd"),
   589 => (x"e2",x"c2",x"87",x"ed"),
   590 => (x"e1",x"c2",x"48",x"c3"),
   591 => (x"c2",x"78",x"bf",x"f7"),
   592 => (x"c2",x"48",x"c7",x"e2"),
   593 => (x"78",x"bf",x"fb",x"e1"),
   594 => (x"bf",x"e2",x"dd",x"c2"),
   595 => (x"c2",x"87",x"c9",x"02"),
   596 => (x"49",x"bf",x"da",x"dd"),
   597 => (x"87",x"c7",x"31",x"c4"),
   598 => (x"bf",x"ff",x"e1",x"c2"),
   599 => (x"c2",x"31",x"c4",x"49"),
   600 => (x"f6",x"59",x"ea",x"dd"),
   601 => (x"5e",x"0e",x"87",x"e9"),
   602 => (x"71",x"0e",x"5c",x"5b"),
   603 => (x"72",x"4b",x"c0",x"4a"),
   604 => (x"e1",x"c0",x"02",x"9a"),
   605 => (x"49",x"a2",x"da",x"87"),
   606 => (x"c2",x"4b",x"69",x"9f"),
   607 => (x"02",x"bf",x"e2",x"dd"),
   608 => (x"a2",x"d4",x"87",x"cf"),
   609 => (x"49",x"69",x"9f",x"49"),
   610 => (x"ff",x"ff",x"c0",x"4c"),
   611 => (x"c2",x"34",x"d0",x"9c"),
   612 => (x"74",x"4c",x"c0",x"87"),
   613 => (x"49",x"73",x"b3",x"49"),
   614 => (x"f5",x"87",x"ed",x"fd"),
   615 => (x"5e",x"0e",x"87",x"ef"),
   616 => (x"0e",x"5d",x"5c",x"5b"),
   617 => (x"4a",x"71",x"86",x"f4"),
   618 => (x"9a",x"72",x"7e",x"c0"),
   619 => (x"c2",x"87",x"d8",x"02"),
   620 => (x"c0",x"48",x"d6",x"d5"),
   621 => (x"ce",x"d5",x"c2",x"78"),
   622 => (x"c7",x"e2",x"c2",x"48"),
   623 => (x"d5",x"c2",x"78",x"bf"),
   624 => (x"e2",x"c2",x"48",x"d2"),
   625 => (x"c2",x"78",x"bf",x"c3"),
   626 => (x"c0",x"48",x"f7",x"dd"),
   627 => (x"e6",x"dd",x"c2",x"50"),
   628 => (x"d5",x"c2",x"49",x"bf"),
   629 => (x"71",x"4a",x"bf",x"d6"),
   630 => (x"c9",x"c4",x"03",x"aa"),
   631 => (x"cf",x"49",x"72",x"87"),
   632 => (x"e9",x"c0",x"05",x"99"),
   633 => (x"f9",x"ed",x"c0",x"87"),
   634 => (x"ce",x"d5",x"c2",x"48"),
   635 => (x"d5",x"c2",x"78",x"bf"),
   636 => (x"d5",x"c2",x"1e",x"da"),
   637 => (x"c2",x"49",x"bf",x"ce"),
   638 => (x"c1",x"48",x"ce",x"d5"),
   639 => (x"e6",x"71",x"78",x"a1"),
   640 => (x"86",x"c4",x"87",x"cb"),
   641 => (x"48",x"f5",x"ed",x"c0"),
   642 => (x"78",x"da",x"d5",x"c2"),
   643 => (x"ed",x"c0",x"87",x"cc"),
   644 => (x"c0",x"48",x"bf",x"f5"),
   645 => (x"ed",x"c0",x"80",x"e0"),
   646 => (x"d5",x"c2",x"58",x"f9"),
   647 => (x"c1",x"48",x"bf",x"d6"),
   648 => (x"da",x"d5",x"c2",x"80"),
   649 => (x"0b",x"75",x"27",x"58"),
   650 => (x"97",x"bf",x"00",x"00"),
   651 => (x"02",x"9d",x"4d",x"bf"),
   652 => (x"c3",x"87",x"e3",x"c2"),
   653 => (x"c2",x"02",x"ad",x"e5"),
   654 => (x"ed",x"c0",x"87",x"dc"),
   655 => (x"cb",x"4b",x"bf",x"f5"),
   656 => (x"4c",x"11",x"49",x"a3"),
   657 => (x"c1",x"05",x"ac",x"cf"),
   658 => (x"49",x"75",x"87",x"d2"),
   659 => (x"89",x"c1",x"99",x"df"),
   660 => (x"dd",x"c2",x"91",x"cd"),
   661 => (x"a3",x"c1",x"81",x"ea"),
   662 => (x"c3",x"51",x"12",x"4a"),
   663 => (x"51",x"12",x"4a",x"a3"),
   664 => (x"12",x"4a",x"a3",x"c5"),
   665 => (x"4a",x"a3",x"c7",x"51"),
   666 => (x"a3",x"c9",x"51",x"12"),
   667 => (x"ce",x"51",x"12",x"4a"),
   668 => (x"51",x"12",x"4a",x"a3"),
   669 => (x"12",x"4a",x"a3",x"d0"),
   670 => (x"4a",x"a3",x"d2",x"51"),
   671 => (x"a3",x"d4",x"51",x"12"),
   672 => (x"d6",x"51",x"12",x"4a"),
   673 => (x"51",x"12",x"4a",x"a3"),
   674 => (x"12",x"4a",x"a3",x"d8"),
   675 => (x"4a",x"a3",x"dc",x"51"),
   676 => (x"a3",x"de",x"51",x"12"),
   677 => (x"c1",x"51",x"12",x"4a"),
   678 => (x"87",x"fa",x"c0",x"7e"),
   679 => (x"99",x"c8",x"49",x"74"),
   680 => (x"87",x"eb",x"c0",x"05"),
   681 => (x"99",x"d0",x"49",x"74"),
   682 => (x"dc",x"87",x"d1",x"05"),
   683 => (x"cb",x"c0",x"02",x"66"),
   684 => (x"dc",x"49",x"73",x"87"),
   685 => (x"98",x"70",x"0f",x"66"),
   686 => (x"87",x"d3",x"c0",x"02"),
   687 => (x"c6",x"c0",x"05",x"6e"),
   688 => (x"ea",x"dd",x"c2",x"87"),
   689 => (x"c0",x"50",x"c0",x"48"),
   690 => (x"48",x"bf",x"f5",x"ed"),
   691 => (x"c2",x"87",x"e1",x"c2"),
   692 => (x"c0",x"48",x"f7",x"dd"),
   693 => (x"dd",x"c2",x"7e",x"50"),
   694 => (x"c2",x"49",x"bf",x"e6"),
   695 => (x"4a",x"bf",x"d6",x"d5"),
   696 => (x"fb",x"04",x"aa",x"71"),
   697 => (x"e2",x"c2",x"87",x"f7"),
   698 => (x"c0",x"05",x"bf",x"c7"),
   699 => (x"dd",x"c2",x"87",x"c8"),
   700 => (x"c1",x"02",x"bf",x"e2"),
   701 => (x"d5",x"c2",x"87",x"f8"),
   702 => (x"f0",x"49",x"bf",x"d2"),
   703 => (x"49",x"70",x"87",x"d5"),
   704 => (x"59",x"d6",x"d5",x"c2"),
   705 => (x"c2",x"48",x"a6",x"c4"),
   706 => (x"78",x"bf",x"d2",x"d5"),
   707 => (x"bf",x"e2",x"dd",x"c2"),
   708 => (x"87",x"d8",x"c0",x"02"),
   709 => (x"cf",x"49",x"66",x"c4"),
   710 => (x"f8",x"ff",x"ff",x"ff"),
   711 => (x"c0",x"02",x"a9",x"99"),
   712 => (x"4c",x"c0",x"87",x"c5"),
   713 => (x"c1",x"87",x"e1",x"c0"),
   714 => (x"87",x"dc",x"c0",x"4c"),
   715 => (x"cf",x"49",x"66",x"c4"),
   716 => (x"a9",x"99",x"f8",x"ff"),
   717 => (x"87",x"c8",x"c0",x"02"),
   718 => (x"c0",x"48",x"a6",x"c8"),
   719 => (x"87",x"c5",x"c0",x"78"),
   720 => (x"c1",x"48",x"a6",x"c8"),
   721 => (x"4c",x"66",x"c8",x"78"),
   722 => (x"c0",x"05",x"9c",x"74"),
   723 => (x"66",x"c4",x"87",x"e0"),
   724 => (x"c2",x"89",x"c2",x"49"),
   725 => (x"4a",x"bf",x"da",x"dd"),
   726 => (x"f3",x"e1",x"c2",x"91"),
   727 => (x"d5",x"c2",x"4a",x"bf"),
   728 => (x"a1",x"72",x"48",x"ce"),
   729 => (x"d6",x"d5",x"c2",x"78"),
   730 => (x"f9",x"78",x"c0",x"48"),
   731 => (x"48",x"c0",x"87",x"df"),
   732 => (x"d6",x"ee",x"8e",x"f4"),
   733 => (x"00",x"00",x"00",x"87"),
   734 => (x"ff",x"ff",x"ff",x"00"),
   735 => (x"00",x"0b",x"85",x"ff"),
   736 => (x"00",x"0b",x"8e",x"00"),
   737 => (x"54",x"41",x"46",x"00"),
   738 => (x"20",x"20",x"32",x"33"),
   739 => (x"41",x"46",x"00",x"20"),
   740 => (x"20",x"36",x"31",x"54"),
   741 => (x"1e",x"00",x"20",x"20"),
   742 => (x"c3",x"48",x"d4",x"ff"),
   743 => (x"48",x"68",x"78",x"ff"),
   744 => (x"ff",x"1e",x"4f",x"26"),
   745 => (x"ff",x"c3",x"48",x"d4"),
   746 => (x"48",x"d0",x"ff",x"78"),
   747 => (x"ff",x"78",x"e1",x"c0"),
   748 => (x"78",x"d4",x"48",x"d4"),
   749 => (x"48",x"cb",x"e2",x"c2"),
   750 => (x"50",x"bf",x"d4",x"ff"),
   751 => (x"ff",x"1e",x"4f",x"26"),
   752 => (x"e0",x"c0",x"48",x"d0"),
   753 => (x"1e",x"4f",x"26",x"78"),
   754 => (x"70",x"87",x"cc",x"ff"),
   755 => (x"c6",x"02",x"99",x"49"),
   756 => (x"a9",x"fb",x"c0",x"87"),
   757 => (x"71",x"87",x"f1",x"05"),
   758 => (x"0e",x"4f",x"26",x"48"),
   759 => (x"0e",x"5c",x"5b",x"5e"),
   760 => (x"4c",x"c0",x"4b",x"71"),
   761 => (x"70",x"87",x"f0",x"fe"),
   762 => (x"c0",x"02",x"99",x"49"),
   763 => (x"ec",x"c0",x"87",x"f9"),
   764 => (x"f2",x"c0",x"02",x"a9"),
   765 => (x"a9",x"fb",x"c0",x"87"),
   766 => (x"87",x"eb",x"c0",x"02"),
   767 => (x"ac",x"b7",x"66",x"cc"),
   768 => (x"d0",x"87",x"c7",x"03"),
   769 => (x"87",x"c2",x"02",x"66"),
   770 => (x"99",x"71",x"53",x"71"),
   771 => (x"c1",x"87",x"c2",x"02"),
   772 => (x"87",x"c3",x"fe",x"84"),
   773 => (x"02",x"99",x"49",x"70"),
   774 => (x"ec",x"c0",x"87",x"cd"),
   775 => (x"87",x"c7",x"02",x"a9"),
   776 => (x"05",x"a9",x"fb",x"c0"),
   777 => (x"d0",x"87",x"d5",x"ff"),
   778 => (x"87",x"c3",x"02",x"66"),
   779 => (x"c0",x"7b",x"97",x"c0"),
   780 => (x"c4",x"05",x"a9",x"ec"),
   781 => (x"c5",x"4a",x"74",x"87"),
   782 => (x"c0",x"4a",x"74",x"87"),
   783 => (x"48",x"72",x"8a",x"0a"),
   784 => (x"4d",x"26",x"87",x"c2"),
   785 => (x"4b",x"26",x"4c",x"26"),
   786 => (x"fd",x"1e",x"4f",x"26"),
   787 => (x"49",x"70",x"87",x"c9"),
   788 => (x"a9",x"b7",x"f0",x"c0"),
   789 => (x"c0",x"87",x"ca",x"04"),
   790 => (x"01",x"a9",x"b7",x"f9"),
   791 => (x"f0",x"c0",x"87",x"c3"),
   792 => (x"b7",x"c1",x"c1",x"89"),
   793 => (x"87",x"ca",x"04",x"a9"),
   794 => (x"a9",x"b7",x"da",x"c1"),
   795 => (x"c0",x"87",x"c3",x"01"),
   796 => (x"48",x"71",x"89",x"f7"),
   797 => (x"5e",x"0e",x"4f",x"26"),
   798 => (x"71",x"0e",x"5c",x"5b"),
   799 => (x"4c",x"d4",x"ff",x"4a"),
   800 => (x"e9",x"c0",x"49",x"72"),
   801 => (x"9b",x"4b",x"70",x"87"),
   802 => (x"c1",x"87",x"c2",x"02"),
   803 => (x"48",x"d0",x"ff",x"8b"),
   804 => (x"d5",x"c1",x"78",x"c5"),
   805 => (x"c6",x"49",x"73",x"7c"),
   806 => (x"df",x"dc",x"c1",x"31"),
   807 => (x"48",x"4a",x"bf",x"97"),
   808 => (x"7c",x"70",x"b0",x"71"),
   809 => (x"c4",x"48",x"d0",x"ff"),
   810 => (x"fe",x"48",x"73",x"78"),
   811 => (x"5e",x"0e",x"87",x"d6"),
   812 => (x"0e",x"5d",x"5c",x"5b"),
   813 => (x"4c",x"71",x"86",x"f8"),
   814 => (x"e5",x"fb",x"7e",x"c0"),
   815 => (x"c0",x"4b",x"c0",x"87"),
   816 => (x"bf",x"97",x"db",x"f5"),
   817 => (x"04",x"a9",x"c0",x"49"),
   818 => (x"fa",x"fb",x"87",x"cf"),
   819 => (x"c0",x"83",x"c1",x"87"),
   820 => (x"bf",x"97",x"db",x"f5"),
   821 => (x"f1",x"06",x"ab",x"49"),
   822 => (x"db",x"f5",x"c0",x"87"),
   823 => (x"cf",x"02",x"bf",x"97"),
   824 => (x"87",x"f3",x"fa",x"87"),
   825 => (x"02",x"99",x"49",x"70"),
   826 => (x"ec",x"c0",x"87",x"c6"),
   827 => (x"87",x"f1",x"05",x"a9"),
   828 => (x"e2",x"fa",x"4b",x"c0"),
   829 => (x"fa",x"4d",x"70",x"87"),
   830 => (x"a6",x"c8",x"87",x"dd"),
   831 => (x"87",x"d7",x"fa",x"58"),
   832 => (x"83",x"c1",x"4a",x"70"),
   833 => (x"97",x"49",x"a4",x"c8"),
   834 => (x"02",x"ad",x"49",x"69"),
   835 => (x"ff",x"c0",x"87",x"c7"),
   836 => (x"e7",x"c0",x"05",x"ad"),
   837 => (x"49",x"a4",x"c9",x"87"),
   838 => (x"c4",x"49",x"69",x"97"),
   839 => (x"c7",x"02",x"a9",x"66"),
   840 => (x"ff",x"c0",x"48",x"87"),
   841 => (x"87",x"d4",x"05",x"a8"),
   842 => (x"97",x"49",x"a4",x"ca"),
   843 => (x"02",x"aa",x"49",x"69"),
   844 => (x"ff",x"c0",x"87",x"c6"),
   845 => (x"87",x"c4",x"05",x"aa"),
   846 => (x"87",x"d0",x"7e",x"c1"),
   847 => (x"02",x"ad",x"ec",x"c0"),
   848 => (x"fb",x"c0",x"87",x"c6"),
   849 => (x"87",x"c4",x"05",x"ad"),
   850 => (x"7e",x"c1",x"4b",x"c0"),
   851 => (x"e1",x"fe",x"02",x"6e"),
   852 => (x"87",x"ea",x"f9",x"87"),
   853 => (x"8e",x"f8",x"48",x"73"),
   854 => (x"00",x"87",x"e7",x"fb"),
   855 => (x"5c",x"5b",x"5e",x"0e"),
   856 => (x"71",x"1e",x"0e",x"5d"),
   857 => (x"4b",x"d4",x"ff",x"4d"),
   858 => (x"e2",x"c2",x"1e",x"75"),
   859 => (x"f3",x"e9",x"49",x"d0"),
   860 => (x"70",x"86",x"c4",x"87"),
   861 => (x"d5",x"c3",x"02",x"98"),
   862 => (x"d8",x"e2",x"c2",x"87"),
   863 => (x"49",x"75",x"4c",x"bf"),
   864 => (x"ff",x"87",x"f3",x"fb"),
   865 => (x"78",x"c5",x"48",x"d0"),
   866 => (x"c0",x"7b",x"d6",x"c1"),
   867 => (x"49",x"a2",x"75",x"4a"),
   868 => (x"82",x"c1",x"7b",x"11"),
   869 => (x"04",x"aa",x"b7",x"cb"),
   870 => (x"4a",x"cc",x"87",x"f3"),
   871 => (x"c1",x"7b",x"ff",x"c3"),
   872 => (x"b7",x"e0",x"c0",x"82"),
   873 => (x"87",x"f4",x"04",x"aa"),
   874 => (x"c4",x"48",x"d0",x"ff"),
   875 => (x"7b",x"ff",x"c3",x"78"),
   876 => (x"d3",x"c1",x"78",x"c5"),
   877 => (x"c4",x"7b",x"c1",x"7b"),
   878 => (x"02",x"9c",x"74",x"78"),
   879 => (x"c2",x"87",x"ff",x"c1"),
   880 => (x"c8",x"7e",x"da",x"d5"),
   881 => (x"c0",x"8c",x"4d",x"c0"),
   882 => (x"c6",x"03",x"ac",x"b7"),
   883 => (x"a4",x"c0",x"c8",x"87"),
   884 => (x"c8",x"4c",x"c0",x"4d"),
   885 => (x"dc",x"05",x"ad",x"c0"),
   886 => (x"cb",x"e2",x"c2",x"87"),
   887 => (x"d0",x"49",x"bf",x"97"),
   888 => (x"87",x"d1",x"02",x"99"),
   889 => (x"e2",x"c2",x"1e",x"c0"),
   890 => (x"cc",x"eb",x"49",x"d0"),
   891 => (x"70",x"86",x"c4",x"87"),
   892 => (x"ee",x"c0",x"4a",x"49"),
   893 => (x"da",x"d5",x"c2",x"87"),
   894 => (x"d0",x"e2",x"c2",x"1e"),
   895 => (x"87",x"f9",x"ea",x"49"),
   896 => (x"49",x"70",x"86",x"c4"),
   897 => (x"48",x"d0",x"ff",x"4a"),
   898 => (x"c1",x"78",x"c5",x"c8"),
   899 => (x"97",x"6e",x"7b",x"d4"),
   900 => (x"48",x"6e",x"7b",x"bf"),
   901 => (x"7e",x"70",x"80",x"c1"),
   902 => (x"ff",x"05",x"8d",x"c1"),
   903 => (x"d0",x"ff",x"87",x"f0"),
   904 => (x"72",x"78",x"c4",x"48"),
   905 => (x"87",x"c5",x"05",x"9a"),
   906 => (x"e3",x"c0",x"48",x"c0"),
   907 => (x"c2",x"1e",x"c1",x"87"),
   908 => (x"e8",x"49",x"d0",x"e2"),
   909 => (x"86",x"c4",x"87",x"e9"),
   910 => (x"fe",x"05",x"9c",x"74"),
   911 => (x"d0",x"ff",x"87",x"c1"),
   912 => (x"c1",x"78",x"c5",x"48"),
   913 => (x"7b",x"c0",x"7b",x"d3"),
   914 => (x"48",x"c1",x"78",x"c4"),
   915 => (x"48",x"c0",x"87",x"c2"),
   916 => (x"26",x"4d",x"26",x"26"),
   917 => (x"26",x"4b",x"26",x"4c"),
   918 => (x"5b",x"5e",x"0e",x"4f"),
   919 => (x"1e",x"0e",x"5d",x"5c"),
   920 => (x"4c",x"c0",x"4b",x"71"),
   921 => (x"c0",x"04",x"ab",x"4d"),
   922 => (x"f2",x"c0",x"87",x"e8"),
   923 => (x"9d",x"75",x"1e",x"ee"),
   924 => (x"c0",x"87",x"c4",x"02"),
   925 => (x"c1",x"87",x"c2",x"4a"),
   926 => (x"ec",x"49",x"72",x"4a"),
   927 => (x"86",x"c4",x"87",x"e0"),
   928 => (x"84",x"c1",x"7e",x"70"),
   929 => (x"87",x"c2",x"05",x"6e"),
   930 => (x"85",x"c1",x"4c",x"73"),
   931 => (x"ff",x"06",x"ac",x"73"),
   932 => (x"48",x"6e",x"87",x"d8"),
   933 => (x"87",x"f9",x"fe",x"26"),
   934 => (x"c4",x"4a",x"71",x"1e"),
   935 => (x"87",x"c5",x"05",x"66"),
   936 => (x"f7",x"fa",x"49",x"72"),
   937 => (x"0e",x"4f",x"26",x"87"),
   938 => (x"5d",x"5c",x"5b",x"5e"),
   939 => (x"4c",x"71",x"1e",x"0e"),
   940 => (x"c2",x"91",x"de",x"49"),
   941 => (x"71",x"4d",x"f8",x"e2"),
   942 => (x"02",x"6d",x"97",x"85"),
   943 => (x"c2",x"87",x"dc",x"c1"),
   944 => (x"4a",x"bf",x"e4",x"e2"),
   945 => (x"49",x"72",x"82",x"74"),
   946 => (x"70",x"87",x"ce",x"fe"),
   947 => (x"c0",x"02",x"6e",x"7e"),
   948 => (x"e2",x"c2",x"87",x"f2"),
   949 => (x"4a",x"6e",x"4b",x"ec"),
   950 => (x"c7",x"ff",x"49",x"cb"),
   951 => (x"4b",x"74",x"87",x"ca"),
   952 => (x"dc",x"c1",x"93",x"cb"),
   953 => (x"83",x"c4",x"83",x"ef"),
   954 => (x"7b",x"df",x"fc",x"c0"),
   955 => (x"c0",x"c1",x"49",x"74"),
   956 => (x"7b",x"75",x"87",x"f4"),
   957 => (x"97",x"e0",x"dc",x"c1"),
   958 => (x"c2",x"1e",x"49",x"bf"),
   959 => (x"fe",x"49",x"ec",x"e2"),
   960 => (x"86",x"c4",x"87",x"d6"),
   961 => (x"c0",x"c1",x"49",x"74"),
   962 => (x"49",x"c0",x"87",x"dc"),
   963 => (x"87",x"fb",x"c1",x"c1"),
   964 => (x"48",x"cc",x"e2",x"c2"),
   965 => (x"49",x"c1",x"78",x"c0"),
   966 => (x"26",x"87",x"c0",x"dd"),
   967 => (x"4c",x"87",x"f2",x"fc"),
   968 => (x"69",x"64",x"61",x"6f"),
   969 => (x"2e",x"2e",x"67",x"6e"),
   970 => (x"5e",x"0e",x"00",x"2e"),
   971 => (x"71",x"0e",x"5c",x"5b"),
   972 => (x"e2",x"c2",x"4a",x"4b"),
   973 => (x"72",x"82",x"bf",x"e4"),
   974 => (x"87",x"dd",x"fc",x"49"),
   975 => (x"02",x"9c",x"4c",x"70"),
   976 => (x"e8",x"49",x"87",x"c4"),
   977 => (x"e2",x"c2",x"87",x"e0"),
   978 => (x"78",x"c0",x"48",x"e4"),
   979 => (x"ca",x"dc",x"49",x"c1"),
   980 => (x"87",x"ff",x"fb",x"87"),
   981 => (x"5c",x"5b",x"5e",x"0e"),
   982 => (x"86",x"f4",x"0e",x"5d"),
   983 => (x"4d",x"da",x"d5",x"c2"),
   984 => (x"a6",x"c4",x"4c",x"c0"),
   985 => (x"c2",x"78",x"c0",x"48"),
   986 => (x"49",x"bf",x"e4",x"e2"),
   987 => (x"c1",x"06",x"a9",x"c0"),
   988 => (x"d5",x"c2",x"87",x"c1"),
   989 => (x"02",x"98",x"48",x"da"),
   990 => (x"c0",x"87",x"f8",x"c0"),
   991 => (x"c8",x"1e",x"ee",x"f2"),
   992 => (x"87",x"c7",x"02",x"66"),
   993 => (x"c0",x"48",x"a6",x"c4"),
   994 => (x"c4",x"87",x"c5",x"78"),
   995 => (x"78",x"c1",x"48",x"a6"),
   996 => (x"e8",x"49",x"66",x"c4"),
   997 => (x"86",x"c4",x"87",x"c8"),
   998 => (x"84",x"c1",x"4d",x"70"),
   999 => (x"c1",x"48",x"66",x"c4"),
  1000 => (x"58",x"a6",x"c8",x"80"),
  1001 => (x"bf",x"e4",x"e2",x"c2"),
  1002 => (x"c6",x"03",x"ac",x"49"),
  1003 => (x"05",x"9d",x"75",x"87"),
  1004 => (x"c0",x"87",x"c8",x"ff"),
  1005 => (x"02",x"9d",x"75",x"4c"),
  1006 => (x"c0",x"87",x"e0",x"c3"),
  1007 => (x"c8",x"1e",x"ee",x"f2"),
  1008 => (x"87",x"c7",x"02",x"66"),
  1009 => (x"c0",x"48",x"a6",x"cc"),
  1010 => (x"cc",x"87",x"c5",x"78"),
  1011 => (x"78",x"c1",x"48",x"a6"),
  1012 => (x"e7",x"49",x"66",x"cc"),
  1013 => (x"86",x"c4",x"87",x"c8"),
  1014 => (x"02",x"6e",x"7e",x"70"),
  1015 => (x"6e",x"87",x"e9",x"c2"),
  1016 => (x"97",x"81",x"cb",x"49"),
  1017 => (x"99",x"d0",x"49",x"69"),
  1018 => (x"87",x"d6",x"c1",x"02"),
  1019 => (x"4a",x"ea",x"fc",x"c0"),
  1020 => (x"91",x"cb",x"49",x"74"),
  1021 => (x"81",x"ef",x"dc",x"c1"),
  1022 => (x"81",x"c8",x"79",x"72"),
  1023 => (x"74",x"51",x"ff",x"c3"),
  1024 => (x"c2",x"91",x"de",x"49"),
  1025 => (x"71",x"4d",x"f8",x"e2"),
  1026 => (x"97",x"c1",x"c2",x"85"),
  1027 => (x"49",x"a5",x"c1",x"7d"),
  1028 => (x"c2",x"51",x"e0",x"c0"),
  1029 => (x"bf",x"97",x"ea",x"dd"),
  1030 => (x"c1",x"87",x"d2",x"02"),
  1031 => (x"4b",x"a5",x"c2",x"84"),
  1032 => (x"4a",x"ea",x"dd",x"c2"),
  1033 => (x"c1",x"ff",x"49",x"db"),
  1034 => (x"db",x"c1",x"87",x"fe"),
  1035 => (x"49",x"a5",x"cd",x"87"),
  1036 => (x"84",x"c1",x"51",x"c0"),
  1037 => (x"6e",x"4b",x"a5",x"c2"),
  1038 => (x"ff",x"49",x"cb",x"4a"),
  1039 => (x"c1",x"87",x"e9",x"c1"),
  1040 => (x"fa",x"c0",x"87",x"c6"),
  1041 => (x"49",x"74",x"4a",x"e7"),
  1042 => (x"dc",x"c1",x"91",x"cb"),
  1043 => (x"79",x"72",x"81",x"ef"),
  1044 => (x"97",x"ea",x"dd",x"c2"),
  1045 => (x"87",x"d8",x"02",x"bf"),
  1046 => (x"91",x"de",x"49",x"74"),
  1047 => (x"e2",x"c2",x"84",x"c1"),
  1048 => (x"83",x"71",x"4b",x"f8"),
  1049 => (x"4a",x"ea",x"dd",x"c2"),
  1050 => (x"c0",x"ff",x"49",x"dd"),
  1051 => (x"87",x"d8",x"87",x"fa"),
  1052 => (x"93",x"de",x"4b",x"74"),
  1053 => (x"83",x"f8",x"e2",x"c2"),
  1054 => (x"c0",x"49",x"a3",x"cb"),
  1055 => (x"73",x"84",x"c1",x"51"),
  1056 => (x"49",x"cb",x"4a",x"6e"),
  1057 => (x"87",x"e0",x"c0",x"ff"),
  1058 => (x"c1",x"48",x"66",x"c4"),
  1059 => (x"58",x"a6",x"c8",x"80"),
  1060 => (x"c0",x"03",x"ac",x"c7"),
  1061 => (x"05",x"6e",x"87",x"c5"),
  1062 => (x"74",x"87",x"e0",x"fc"),
  1063 => (x"f6",x"8e",x"f4",x"48"),
  1064 => (x"73",x"1e",x"87",x"ef"),
  1065 => (x"49",x"4b",x"71",x"1e"),
  1066 => (x"dc",x"c1",x"91",x"cb"),
  1067 => (x"a1",x"c8",x"81",x"ef"),
  1068 => (x"df",x"dc",x"c1",x"4a"),
  1069 => (x"c9",x"50",x"12",x"48"),
  1070 => (x"f5",x"c0",x"4a",x"a1"),
  1071 => (x"50",x"12",x"48",x"db"),
  1072 => (x"dc",x"c1",x"81",x"ca"),
  1073 => (x"50",x"11",x"48",x"e0"),
  1074 => (x"97",x"e0",x"dc",x"c1"),
  1075 => (x"c0",x"1e",x"49",x"bf"),
  1076 => (x"87",x"c4",x"f7",x"49"),
  1077 => (x"48",x"cc",x"e2",x"c2"),
  1078 => (x"49",x"c1",x"78",x"de"),
  1079 => (x"26",x"87",x"fc",x"d5"),
  1080 => (x"1e",x"87",x"f2",x"f5"),
  1081 => (x"cb",x"49",x"4a",x"71"),
  1082 => (x"ef",x"dc",x"c1",x"91"),
  1083 => (x"11",x"81",x"c8",x"81"),
  1084 => (x"d0",x"e2",x"c2",x"48"),
  1085 => (x"e4",x"e2",x"c2",x"58"),
  1086 => (x"c1",x"78",x"c0",x"48"),
  1087 => (x"87",x"db",x"d5",x"49"),
  1088 => (x"c0",x"1e",x"4f",x"26"),
  1089 => (x"c2",x"fa",x"c0",x"49"),
  1090 => (x"1e",x"4f",x"26",x"87"),
  1091 => (x"d2",x"02",x"99",x"71"),
  1092 => (x"c4",x"de",x"c1",x"87"),
  1093 => (x"f7",x"50",x"c0",x"48"),
  1094 => (x"e3",x"c3",x"c1",x"80"),
  1095 => (x"e8",x"dc",x"c1",x"40"),
  1096 => (x"c1",x"87",x"ce",x"78"),
  1097 => (x"c1",x"48",x"c0",x"de"),
  1098 => (x"fc",x"78",x"e1",x"dc"),
  1099 => (x"c2",x"c4",x"c1",x"80"),
  1100 => (x"0e",x"4f",x"26",x"78"),
  1101 => (x"0e",x"5c",x"5b",x"5e"),
  1102 => (x"cb",x"4a",x"4c",x"71"),
  1103 => (x"ef",x"dc",x"c1",x"92"),
  1104 => (x"49",x"a2",x"c8",x"82"),
  1105 => (x"97",x"4b",x"a2",x"c9"),
  1106 => (x"97",x"1e",x"4b",x"6b"),
  1107 => (x"ca",x"1e",x"49",x"69"),
  1108 => (x"c0",x"49",x"12",x"82"),
  1109 => (x"c0",x"87",x"fd",x"e4"),
  1110 => (x"87",x"ff",x"d3",x"49"),
  1111 => (x"f7",x"c0",x"49",x"74"),
  1112 => (x"8e",x"f8",x"87",x"c4"),
  1113 => (x"1e",x"87",x"ec",x"f3"),
  1114 => (x"4b",x"71",x"1e",x"73"),
  1115 => (x"87",x"c3",x"ff",x"49"),
  1116 => (x"fe",x"fe",x"49",x"73"),
  1117 => (x"87",x"dd",x"f3",x"87"),
  1118 => (x"71",x"1e",x"73",x"1e"),
  1119 => (x"4a",x"a3",x"c6",x"4b"),
  1120 => (x"c1",x"87",x"db",x"02"),
  1121 => (x"87",x"d6",x"02",x"8a"),
  1122 => (x"da",x"c1",x"02",x"8a"),
  1123 => (x"c0",x"02",x"8a",x"87"),
  1124 => (x"02",x"8a",x"87",x"fc"),
  1125 => (x"8a",x"87",x"e1",x"c0"),
  1126 => (x"c1",x"87",x"cb",x"02"),
  1127 => (x"49",x"c7",x"87",x"db"),
  1128 => (x"c1",x"87",x"c0",x"fd"),
  1129 => (x"e2",x"c2",x"87",x"de"),
  1130 => (x"c1",x"02",x"bf",x"e4"),
  1131 => (x"c1",x"48",x"87",x"cb"),
  1132 => (x"e8",x"e2",x"c2",x"88"),
  1133 => (x"87",x"c1",x"c1",x"58"),
  1134 => (x"bf",x"e8",x"e2",x"c2"),
  1135 => (x"87",x"f9",x"c0",x"02"),
  1136 => (x"bf",x"e4",x"e2",x"c2"),
  1137 => (x"c2",x"80",x"c1",x"48"),
  1138 => (x"c0",x"58",x"e8",x"e2"),
  1139 => (x"e2",x"c2",x"87",x"eb"),
  1140 => (x"c6",x"49",x"bf",x"e4"),
  1141 => (x"e8",x"e2",x"c2",x"89"),
  1142 => (x"a9",x"b7",x"c0",x"59"),
  1143 => (x"c2",x"87",x"da",x"03"),
  1144 => (x"c0",x"48",x"e4",x"e2"),
  1145 => (x"c2",x"87",x"d2",x"78"),
  1146 => (x"02",x"bf",x"e8",x"e2"),
  1147 => (x"e2",x"c2",x"87",x"cb"),
  1148 => (x"c6",x"48",x"bf",x"e4"),
  1149 => (x"e8",x"e2",x"c2",x"80"),
  1150 => (x"d1",x"49",x"c0",x"58"),
  1151 => (x"49",x"73",x"87",x"dd"),
  1152 => (x"87",x"e2",x"f4",x"c0"),
  1153 => (x"0e",x"87",x"ce",x"f1"),
  1154 => (x"0e",x"5c",x"5b",x"5e"),
  1155 => (x"66",x"cc",x"4c",x"71"),
  1156 => (x"cb",x"4b",x"74",x"1e"),
  1157 => (x"ef",x"dc",x"c1",x"93"),
  1158 => (x"4a",x"a3",x"c4",x"83"),
  1159 => (x"fa",x"fe",x"49",x"6a"),
  1160 => (x"c2",x"c1",x"87",x"d6"),
  1161 => (x"a3",x"c8",x"7b",x"e2"),
  1162 => (x"51",x"66",x"d4",x"49"),
  1163 => (x"d8",x"49",x"a3",x"c9"),
  1164 => (x"a3",x"ca",x"51",x"66"),
  1165 => (x"51",x"66",x"dc",x"49"),
  1166 => (x"87",x"d7",x"f0",x"26"),
  1167 => (x"5c",x"5b",x"5e",x"0e"),
  1168 => (x"d0",x"ff",x"0e",x"5d"),
  1169 => (x"59",x"a6",x"d8",x"86"),
  1170 => (x"c0",x"48",x"a6",x"c4"),
  1171 => (x"c1",x"80",x"c4",x"78"),
  1172 => (x"c4",x"78",x"66",x"c4"),
  1173 => (x"c4",x"78",x"c1",x"80"),
  1174 => (x"c2",x"78",x"c1",x"80"),
  1175 => (x"c1",x"48",x"e8",x"e2"),
  1176 => (x"cc",x"e2",x"c2",x"78"),
  1177 => (x"a8",x"de",x"48",x"bf"),
  1178 => (x"f3",x"87",x"cb",x"05"),
  1179 => (x"49",x"70",x"87",x"e6"),
  1180 => (x"ce",x"59",x"a6",x"c8"),
  1181 => (x"e9",x"e4",x"87",x"ed"),
  1182 => (x"87",x"cb",x"e5",x"87"),
  1183 => (x"70",x"87",x"d8",x"e4"),
  1184 => (x"ac",x"fb",x"c0",x"4c"),
  1185 => (x"87",x"d0",x"c1",x"02"),
  1186 => (x"c1",x"05",x"66",x"d4"),
  1187 => (x"1e",x"c0",x"87",x"c2"),
  1188 => (x"c1",x"1e",x"c1",x"1e"),
  1189 => (x"c0",x"1e",x"d2",x"de"),
  1190 => (x"87",x"eb",x"fd",x"49"),
  1191 => (x"4a",x"66",x"d0",x"c1"),
  1192 => (x"49",x"6a",x"82",x"c4"),
  1193 => (x"51",x"74",x"81",x"c7"),
  1194 => (x"1e",x"d8",x"1e",x"c1"),
  1195 => (x"81",x"c8",x"49",x"6a"),
  1196 => (x"d8",x"87",x"e8",x"e4"),
  1197 => (x"66",x"c4",x"c1",x"86"),
  1198 => (x"01",x"a8",x"c0",x"48"),
  1199 => (x"a6",x"c4",x"87",x"c7"),
  1200 => (x"ce",x"78",x"c1",x"48"),
  1201 => (x"66",x"c4",x"c1",x"87"),
  1202 => (x"cc",x"88",x"c1",x"48"),
  1203 => (x"87",x"c3",x"58",x"a6"),
  1204 => (x"cc",x"87",x"f4",x"e3"),
  1205 => (x"78",x"c2",x"48",x"a6"),
  1206 => (x"cd",x"02",x"9c",x"74"),
  1207 => (x"66",x"c4",x"87",x"c1"),
  1208 => (x"66",x"c8",x"c1",x"48"),
  1209 => (x"f6",x"cc",x"03",x"a8"),
  1210 => (x"48",x"a6",x"d8",x"87"),
  1211 => (x"80",x"c4",x"78",x"c0"),
  1212 => (x"e2",x"e2",x"78",x"c0"),
  1213 => (x"c1",x"4c",x"70",x"87"),
  1214 => (x"c2",x"05",x"ac",x"d0"),
  1215 => (x"66",x"dc",x"87",x"d7"),
  1216 => (x"87",x"c6",x"e5",x"7e"),
  1217 => (x"e0",x"c0",x"49",x"70"),
  1218 => (x"ca",x"e2",x"59",x"a6"),
  1219 => (x"c0",x"4c",x"70",x"87"),
  1220 => (x"c1",x"05",x"ac",x"ec"),
  1221 => (x"66",x"c4",x"87",x"ea"),
  1222 => (x"c1",x"91",x"cb",x"49"),
  1223 => (x"c4",x"81",x"66",x"c0"),
  1224 => (x"4d",x"6a",x"4a",x"a1"),
  1225 => (x"dc",x"4a",x"a1",x"c8"),
  1226 => (x"c3",x"c1",x"52",x"66"),
  1227 => (x"e6",x"e1",x"79",x"e3"),
  1228 => (x"9c",x"4c",x"70",x"87"),
  1229 => (x"c0",x"87",x"d8",x"02"),
  1230 => (x"d2",x"02",x"ac",x"fb"),
  1231 => (x"e1",x"55",x"74",x"87"),
  1232 => (x"4c",x"70",x"87",x"d5"),
  1233 => (x"87",x"c7",x"02",x"9c"),
  1234 => (x"05",x"ac",x"fb",x"c0"),
  1235 => (x"c0",x"87",x"ee",x"ff"),
  1236 => (x"c1",x"c2",x"55",x"e0"),
  1237 => (x"7d",x"97",x"c0",x"55"),
  1238 => (x"6e",x"49",x"66",x"d4"),
  1239 => (x"87",x"db",x"05",x"a9"),
  1240 => (x"c8",x"48",x"66",x"c4"),
  1241 => (x"ca",x"04",x"a8",x"66"),
  1242 => (x"48",x"66",x"c4",x"87"),
  1243 => (x"a6",x"c8",x"80",x"c1"),
  1244 => (x"c8",x"87",x"c8",x"58"),
  1245 => (x"88",x"c1",x"48",x"66"),
  1246 => (x"e0",x"58",x"a6",x"cc"),
  1247 => (x"4c",x"70",x"87",x"d9"),
  1248 => (x"05",x"ac",x"d0",x"c1"),
  1249 => (x"66",x"d0",x"87",x"c8"),
  1250 => (x"d4",x"80",x"c1",x"48"),
  1251 => (x"d0",x"c1",x"58",x"a6"),
  1252 => (x"e9",x"fd",x"02",x"ac"),
  1253 => (x"a6",x"e0",x"c0",x"87"),
  1254 => (x"78",x"66",x"d4",x"48"),
  1255 => (x"c0",x"48",x"66",x"dc"),
  1256 => (x"05",x"a8",x"66",x"e0"),
  1257 => (x"c0",x"87",x"ca",x"c9"),
  1258 => (x"c0",x"48",x"a6",x"e4"),
  1259 => (x"48",x"74",x"7e",x"78"),
  1260 => (x"c0",x"88",x"fb",x"c0"),
  1261 => (x"70",x"58",x"a6",x"ec"),
  1262 => (x"cf",x"c8",x"02",x"98"),
  1263 => (x"88",x"cb",x"48",x"87"),
  1264 => (x"58",x"a6",x"ec",x"c0"),
  1265 => (x"c1",x"02",x"98",x"70"),
  1266 => (x"c9",x"48",x"87",x"d2"),
  1267 => (x"a6",x"ec",x"c0",x"88"),
  1268 => (x"02",x"98",x"70",x"58"),
  1269 => (x"48",x"87",x"db",x"c3"),
  1270 => (x"ec",x"c0",x"88",x"c4"),
  1271 => (x"98",x"70",x"58",x"a6"),
  1272 => (x"48",x"87",x"d0",x"02"),
  1273 => (x"ec",x"c0",x"88",x"c1"),
  1274 => (x"98",x"70",x"58",x"a6"),
  1275 => (x"87",x"c2",x"c3",x"02"),
  1276 => (x"d8",x"87",x"d3",x"c7"),
  1277 => (x"f0",x"c0",x"48",x"a6"),
  1278 => (x"da",x"de",x"ff",x"78"),
  1279 => (x"c0",x"4c",x"70",x"87"),
  1280 => (x"c0",x"02",x"ac",x"ec"),
  1281 => (x"a6",x"dc",x"87",x"c3"),
  1282 => (x"ac",x"ec",x"c0",x"5c"),
  1283 => (x"ff",x"87",x"cd",x"02"),
  1284 => (x"70",x"87",x"c4",x"de"),
  1285 => (x"ac",x"ec",x"c0",x"4c"),
  1286 => (x"87",x"f3",x"ff",x"05"),
  1287 => (x"02",x"ac",x"ec",x"c0"),
  1288 => (x"ff",x"87",x"c4",x"c0"),
  1289 => (x"d8",x"87",x"f0",x"dd"),
  1290 => (x"66",x"d4",x"1e",x"66"),
  1291 => (x"66",x"d4",x"1e",x"49"),
  1292 => (x"de",x"c1",x"1e",x"49"),
  1293 => (x"66",x"d4",x"1e",x"d2"),
  1294 => (x"87",x"cb",x"f7",x"49"),
  1295 => (x"1e",x"ca",x"1e",x"c0"),
  1296 => (x"cb",x"49",x"66",x"dc"),
  1297 => (x"66",x"d8",x"c1",x"91"),
  1298 => (x"48",x"a6",x"d8",x"81"),
  1299 => (x"d8",x"78",x"a1",x"c4"),
  1300 => (x"ff",x"49",x"bf",x"66"),
  1301 => (x"d8",x"87",x"c4",x"de"),
  1302 => (x"a8",x"b7",x"c0",x"86"),
  1303 => (x"87",x"c5",x"c1",x"06"),
  1304 => (x"1e",x"de",x"1e",x"c1"),
  1305 => (x"49",x"bf",x"66",x"c8"),
  1306 => (x"87",x"ef",x"dd",x"ff"),
  1307 => (x"49",x"70",x"86",x"c8"),
  1308 => (x"88",x"08",x"c0",x"48"),
  1309 => (x"c0",x"58",x"a6",x"dc"),
  1310 => (x"c0",x"06",x"a8",x"b7"),
  1311 => (x"66",x"d8",x"87",x"e7"),
  1312 => (x"a8",x"b7",x"dd",x"48"),
  1313 => (x"6e",x"87",x"de",x"03"),
  1314 => (x"66",x"d8",x"49",x"bf"),
  1315 => (x"51",x"e0",x"c0",x"81"),
  1316 => (x"c1",x"49",x"66",x"d8"),
  1317 => (x"81",x"bf",x"6e",x"81"),
  1318 => (x"d8",x"51",x"c1",x"c2"),
  1319 => (x"81",x"c2",x"49",x"66"),
  1320 => (x"c0",x"81",x"bf",x"6e"),
  1321 => (x"48",x"66",x"cc",x"51"),
  1322 => (x"a6",x"d0",x"80",x"c1"),
  1323 => (x"c4",x"7e",x"c1",x"58"),
  1324 => (x"de",x"ff",x"87",x"da"),
  1325 => (x"a6",x"dc",x"87",x"d4"),
  1326 => (x"cd",x"de",x"ff",x"58"),
  1327 => (x"a6",x"ec",x"c0",x"87"),
  1328 => (x"a8",x"ec",x"c0",x"58"),
  1329 => (x"87",x"ca",x"c0",x"05"),
  1330 => (x"48",x"a6",x"e8",x"c0"),
  1331 => (x"c0",x"78",x"66",x"d8"),
  1332 => (x"db",x"ff",x"87",x"c4"),
  1333 => (x"66",x"c4",x"87",x"c1"),
  1334 => (x"c1",x"91",x"cb",x"49"),
  1335 => (x"71",x"48",x"66",x"c0"),
  1336 => (x"6e",x"7e",x"70",x"80"),
  1337 => (x"6e",x"82",x"c8",x"4a"),
  1338 => (x"d8",x"81",x"ca",x"49"),
  1339 => (x"e8",x"c0",x"51",x"66"),
  1340 => (x"81",x"c1",x"49",x"66"),
  1341 => (x"c1",x"89",x"66",x"d8"),
  1342 => (x"70",x"30",x"71",x"48"),
  1343 => (x"71",x"89",x"c1",x"49"),
  1344 => (x"e6",x"c2",x"7a",x"97"),
  1345 => (x"d8",x"49",x"bf",x"d4"),
  1346 => (x"6a",x"97",x"29",x"66"),
  1347 => (x"98",x"71",x"48",x"4a"),
  1348 => (x"58",x"a6",x"f0",x"c0"),
  1349 => (x"81",x"c4",x"49",x"6e"),
  1350 => (x"e0",x"c0",x"4d",x"69"),
  1351 => (x"66",x"dc",x"48",x"66"),
  1352 => (x"c8",x"c0",x"02",x"a8"),
  1353 => (x"48",x"a6",x"d8",x"87"),
  1354 => (x"c5",x"c0",x"78",x"c0"),
  1355 => (x"48",x"a6",x"d8",x"87"),
  1356 => (x"66",x"d8",x"78",x"c1"),
  1357 => (x"1e",x"e0",x"c0",x"1e"),
  1358 => (x"da",x"ff",x"49",x"75"),
  1359 => (x"86",x"c8",x"87",x"dd"),
  1360 => (x"b7",x"c0",x"4c",x"70"),
  1361 => (x"d4",x"c1",x"06",x"ac"),
  1362 => (x"c0",x"85",x"74",x"87"),
  1363 => (x"89",x"74",x"49",x"e0"),
  1364 => (x"d9",x"c1",x"4b",x"75"),
  1365 => (x"fe",x"71",x"4a",x"d8"),
  1366 => (x"c2",x"87",x"cd",x"ed"),
  1367 => (x"66",x"e4",x"c0",x"85"),
  1368 => (x"c0",x"80",x"c1",x"48"),
  1369 => (x"c0",x"58",x"a6",x"e8"),
  1370 => (x"c1",x"49",x"66",x"ec"),
  1371 => (x"02",x"a9",x"70",x"81"),
  1372 => (x"d8",x"87",x"c8",x"c0"),
  1373 => (x"78",x"c0",x"48",x"a6"),
  1374 => (x"d8",x"87",x"c5",x"c0"),
  1375 => (x"78",x"c1",x"48",x"a6"),
  1376 => (x"c2",x"1e",x"66",x"d8"),
  1377 => (x"e0",x"c0",x"49",x"a4"),
  1378 => (x"70",x"88",x"71",x"48"),
  1379 => (x"49",x"75",x"1e",x"49"),
  1380 => (x"87",x"c7",x"d9",x"ff"),
  1381 => (x"b7",x"c0",x"86",x"c8"),
  1382 => (x"c0",x"ff",x"01",x"a8"),
  1383 => (x"66",x"e4",x"c0",x"87"),
  1384 => (x"87",x"d1",x"c0",x"02"),
  1385 => (x"81",x"c9",x"49",x"6e"),
  1386 => (x"51",x"66",x"e4",x"c0"),
  1387 => (x"c4",x"c1",x"48",x"6e"),
  1388 => (x"cc",x"c0",x"78",x"f3"),
  1389 => (x"c9",x"49",x"6e",x"87"),
  1390 => (x"6e",x"51",x"c2",x"81"),
  1391 => (x"e7",x"c5",x"c1",x"48"),
  1392 => (x"c0",x"7e",x"c1",x"78"),
  1393 => (x"d7",x"ff",x"87",x"c6"),
  1394 => (x"4c",x"70",x"87",x"fd"),
  1395 => (x"f5",x"c0",x"02",x"6e"),
  1396 => (x"48",x"66",x"c4",x"87"),
  1397 => (x"04",x"a8",x"66",x"c8"),
  1398 => (x"c4",x"87",x"cb",x"c0"),
  1399 => (x"80",x"c1",x"48",x"66"),
  1400 => (x"c0",x"58",x"a6",x"c8"),
  1401 => (x"66",x"c8",x"87",x"e0"),
  1402 => (x"cc",x"88",x"c1",x"48"),
  1403 => (x"d5",x"c0",x"58",x"a6"),
  1404 => (x"ac",x"c6",x"c1",x"87"),
  1405 => (x"87",x"c8",x"c0",x"05"),
  1406 => (x"c1",x"48",x"66",x"cc"),
  1407 => (x"58",x"a6",x"d0",x"80"),
  1408 => (x"87",x"c3",x"d7",x"ff"),
  1409 => (x"66",x"d0",x"4c",x"70"),
  1410 => (x"d4",x"80",x"c1",x"48"),
  1411 => (x"9c",x"74",x"58",x"a6"),
  1412 => (x"87",x"cb",x"c0",x"02"),
  1413 => (x"c1",x"48",x"66",x"c4"),
  1414 => (x"04",x"a8",x"66",x"c8"),
  1415 => (x"ff",x"87",x"ca",x"f3"),
  1416 => (x"c4",x"87",x"db",x"d6"),
  1417 => (x"a8",x"c7",x"48",x"66"),
  1418 => (x"87",x"e5",x"c0",x"03"),
  1419 => (x"48",x"e8",x"e2",x"c2"),
  1420 => (x"66",x"c4",x"78",x"c0"),
  1421 => (x"c1",x"91",x"cb",x"49"),
  1422 => (x"c4",x"81",x"66",x"c0"),
  1423 => (x"4a",x"6a",x"4a",x"a1"),
  1424 => (x"c4",x"79",x"52",x"c0"),
  1425 => (x"80",x"c1",x"48",x"66"),
  1426 => (x"c7",x"58",x"a6",x"c8"),
  1427 => (x"db",x"ff",x"04",x"a8"),
  1428 => (x"8e",x"d0",x"ff",x"87"),
  1429 => (x"87",x"f9",x"df",x"ff"),
  1430 => (x"1e",x"00",x"20",x"3a"),
  1431 => (x"4b",x"71",x"1e",x"73"),
  1432 => (x"87",x"c6",x"02",x"9b"),
  1433 => (x"48",x"e4",x"e2",x"c2"),
  1434 => (x"1e",x"c7",x"78",x"c0"),
  1435 => (x"bf",x"e4",x"e2",x"c2"),
  1436 => (x"dc",x"c1",x"1e",x"49"),
  1437 => (x"e2",x"c2",x"1e",x"ef"),
  1438 => (x"ee",x"49",x"bf",x"cc"),
  1439 => (x"86",x"cc",x"87",x"fe"),
  1440 => (x"bf",x"cc",x"e2",x"c2"),
  1441 => (x"87",x"c3",x"ea",x"49"),
  1442 => (x"c8",x"02",x"9b",x"73"),
  1443 => (x"ef",x"dc",x"c1",x"87"),
  1444 => (x"e3",x"e3",x"c0",x"49"),
  1445 => (x"fc",x"de",x"ff",x"87"),
  1446 => (x"d4",x"c7",x"1e",x"87"),
  1447 => (x"fe",x"49",x"c1",x"87"),
  1448 => (x"f0",x"fe",x"87",x"f9"),
  1449 => (x"98",x"70",x"87",x"d0"),
  1450 => (x"fe",x"87",x"cd",x"02"),
  1451 => (x"70",x"87",x"e9",x"f7"),
  1452 => (x"87",x"c4",x"02",x"98"),
  1453 => (x"87",x"c2",x"4a",x"c1"),
  1454 => (x"9a",x"72",x"4a",x"c0"),
  1455 => (x"c0",x"87",x"ce",x"05"),
  1456 => (x"ea",x"db",x"c1",x"1e"),
  1457 => (x"fa",x"f0",x"c0",x"49"),
  1458 => (x"fe",x"86",x"c4",x"87"),
  1459 => (x"c1",x"1e",x"c0",x"87"),
  1460 => (x"c0",x"49",x"f5",x"db"),
  1461 => (x"c0",x"87",x"ec",x"f0"),
  1462 => (x"d5",x"f6",x"c0",x"1e"),
  1463 => (x"c0",x"49",x"70",x"87"),
  1464 => (x"c3",x"87",x"e0",x"f0"),
  1465 => (x"8e",x"f8",x"87",x"ca"),
  1466 => (x"44",x"53",x"4f",x"26"),
  1467 => (x"69",x"61",x"66",x"20"),
  1468 => (x"2e",x"64",x"65",x"6c"),
  1469 => (x"6f",x"6f",x"42",x"00"),
  1470 => (x"67",x"6e",x"69",x"74"),
  1471 => (x"00",x"2e",x"2e",x"2e"),
  1472 => (x"d4",x"e7",x"c0",x"1e"),
  1473 => (x"26",x"87",x"fa",x"87"),
  1474 => (x"e2",x"c2",x"1e",x"4f"),
  1475 => (x"78",x"c0",x"48",x"e4"),
  1476 => (x"48",x"cc",x"e2",x"c2"),
  1477 => (x"c0",x"fe",x"78",x"c0"),
  1478 => (x"c0",x"87",x"e5",x"87"),
  1479 => (x"00",x"4f",x"26",x"48"),
  1480 => (x"45",x"20",x"80",x"00"),
  1481 => (x"00",x"74",x"69",x"78"),
  1482 => (x"61",x"42",x"20",x"80"),
  1483 => (x"e3",x"00",x"6b",x"63"),
  1484 => (x"b8",x"00",x"00",x"10"),
  1485 => (x"00",x"00",x"00",x"28"),
  1486 => (x"10",x"e3",x"00",x"00"),
  1487 => (x"28",x"d6",x"00",x"00"),
  1488 => (x"00",x"00",x"00",x"00"),
  1489 => (x"00",x"10",x"e3",x"00"),
  1490 => (x"00",x"28",x"f4",x"00"),
  1491 => (x"00",x"00",x"00",x"00"),
  1492 => (x"00",x"00",x"10",x"e3"),
  1493 => (x"00",x"00",x"29",x"12"),
  1494 => (x"e3",x"00",x"00",x"00"),
  1495 => (x"30",x"00",x"00",x"10"),
  1496 => (x"00",x"00",x"00",x"29"),
  1497 => (x"10",x"e3",x"00",x"00"),
  1498 => (x"29",x"4e",x"00",x"00"),
  1499 => (x"00",x"00",x"00",x"00"),
  1500 => (x"00",x"10",x"e3",x"00"),
  1501 => (x"00",x"29",x"6c",x"00"),
  1502 => (x"00",x"00",x"00",x"00"),
  1503 => (x"00",x"00",x"10",x"e3"),
  1504 => (x"00",x"00",x"00",x"00"),
  1505 => (x"78",x"00",x"00",x"00"),
  1506 => (x"00",x"00",x"00",x"11"),
  1507 => (x"00",x"00",x"00",x"00"),
  1508 => (x"6f",x"4c",x"00",x"00"),
  1509 => (x"2a",x"20",x"64",x"61"),
  1510 => (x"fe",x"1e",x"00",x"2e"),
  1511 => (x"78",x"c0",x"48",x"f0"),
  1512 => (x"09",x"79",x"09",x"cd"),
  1513 => (x"1e",x"1e",x"4f",x"26"),
  1514 => (x"7e",x"bf",x"f0",x"fe"),
  1515 => (x"4f",x"26",x"26",x"48"),
  1516 => (x"48",x"f0",x"fe",x"1e"),
  1517 => (x"4f",x"26",x"78",x"c1"),
  1518 => (x"48",x"f0",x"fe",x"1e"),
  1519 => (x"4f",x"26",x"78",x"c0"),
  1520 => (x"c0",x"4a",x"71",x"1e"),
  1521 => (x"4f",x"26",x"52",x"52"),
  1522 => (x"5c",x"5b",x"5e",x"0e"),
  1523 => (x"86",x"f4",x"0e",x"5d"),
  1524 => (x"6d",x"97",x"4d",x"71"),
  1525 => (x"4c",x"a5",x"c1",x"7e"),
  1526 => (x"c8",x"48",x"6c",x"97"),
  1527 => (x"48",x"6e",x"58",x"a6"),
  1528 => (x"05",x"a8",x"66",x"c4"),
  1529 => (x"48",x"ff",x"87",x"c5"),
  1530 => (x"ff",x"87",x"e6",x"c0"),
  1531 => (x"a5",x"c2",x"87",x"ca"),
  1532 => (x"4b",x"6c",x"97",x"49"),
  1533 => (x"97",x"4b",x"a3",x"71"),
  1534 => (x"6c",x"97",x"4b",x"6b"),
  1535 => (x"c1",x"48",x"6e",x"7e"),
  1536 => (x"58",x"a6",x"c8",x"80"),
  1537 => (x"a6",x"cc",x"98",x"c7"),
  1538 => (x"7c",x"97",x"70",x"58"),
  1539 => (x"73",x"87",x"e1",x"fe"),
  1540 => (x"26",x"8e",x"f4",x"48"),
  1541 => (x"26",x"4c",x"26",x"4d"),
  1542 => (x"0e",x"4f",x"26",x"4b"),
  1543 => (x"0e",x"5c",x"5b",x"5e"),
  1544 => (x"4c",x"71",x"86",x"f4"),
  1545 => (x"c3",x"4a",x"66",x"d8"),
  1546 => (x"a4",x"c2",x"9a",x"ff"),
  1547 => (x"49",x"6c",x"97",x"4b"),
  1548 => (x"72",x"49",x"a1",x"73"),
  1549 => (x"7e",x"6c",x"97",x"51"),
  1550 => (x"80",x"c1",x"48",x"6e"),
  1551 => (x"c7",x"58",x"a6",x"c8"),
  1552 => (x"58",x"a6",x"cc",x"98"),
  1553 => (x"8e",x"f4",x"54",x"70"),
  1554 => (x"1e",x"87",x"ca",x"ff"),
  1555 => (x"87",x"e8",x"fd",x"1e"),
  1556 => (x"49",x"4a",x"bf",x"e0"),
  1557 => (x"99",x"c0",x"e0",x"c0"),
  1558 => (x"72",x"87",x"cb",x"02"),
  1559 => (x"ca",x"e6",x"c2",x"1e"),
  1560 => (x"87",x"f7",x"fe",x"49"),
  1561 => (x"fd",x"fc",x"86",x"c4"),
  1562 => (x"fd",x"7e",x"70",x"87"),
  1563 => (x"26",x"26",x"87",x"c2"),
  1564 => (x"e6",x"c2",x"1e",x"4f"),
  1565 => (x"c7",x"fd",x"49",x"ca"),
  1566 => (x"cb",x"e1",x"c1",x"87"),
  1567 => (x"87",x"da",x"fc",x"49"),
  1568 => (x"26",x"87",x"dc",x"c3"),
  1569 => (x"4f",x"26",x"1e",x"4f"),
  1570 => (x"5c",x"5b",x"5e",x"0e"),
  1571 => (x"c2",x"4c",x"71",x"0e"),
  1572 => (x"fc",x"49",x"ca",x"e6"),
  1573 => (x"4a",x"70",x"87",x"f2"),
  1574 => (x"04",x"aa",x"b7",x"c0"),
  1575 => (x"c3",x"87",x"e3",x"c2"),
  1576 => (x"c9",x"05",x"aa",x"e0"),
  1577 => (x"d2",x"e5",x"c1",x"87"),
  1578 => (x"c2",x"78",x"c1",x"48"),
  1579 => (x"f0",x"c3",x"87",x"d4"),
  1580 => (x"87",x"c9",x"05",x"aa"),
  1581 => (x"48",x"ce",x"e5",x"c1"),
  1582 => (x"f5",x"c1",x"78",x"c1"),
  1583 => (x"d2",x"e5",x"c1",x"87"),
  1584 => (x"87",x"c7",x"02",x"bf"),
  1585 => (x"c0",x"c2",x"4b",x"72"),
  1586 => (x"72",x"87",x"c2",x"b3"),
  1587 => (x"05",x"9c",x"74",x"4b"),
  1588 => (x"e5",x"c1",x"87",x"d1"),
  1589 => (x"c1",x"1e",x"bf",x"ce"),
  1590 => (x"1e",x"bf",x"d2",x"e5"),
  1591 => (x"e4",x"fe",x"49",x"72"),
  1592 => (x"c1",x"86",x"c8",x"87"),
  1593 => (x"02",x"bf",x"ce",x"e5"),
  1594 => (x"73",x"87",x"e0",x"c0"),
  1595 => (x"29",x"b7",x"c4",x"49"),
  1596 => (x"ee",x"e6",x"c1",x"91"),
  1597 => (x"cf",x"4a",x"73",x"81"),
  1598 => (x"c1",x"92",x"c2",x"9a"),
  1599 => (x"70",x"30",x"72",x"48"),
  1600 => (x"72",x"ba",x"ff",x"4a"),
  1601 => (x"70",x"98",x"69",x"48"),
  1602 => (x"73",x"87",x"db",x"79"),
  1603 => (x"29",x"b7",x"c4",x"49"),
  1604 => (x"ee",x"e6",x"c1",x"91"),
  1605 => (x"cf",x"4a",x"73",x"81"),
  1606 => (x"c3",x"92",x"c2",x"9a"),
  1607 => (x"70",x"30",x"72",x"48"),
  1608 => (x"b0",x"69",x"48",x"4a"),
  1609 => (x"e5",x"c1",x"79",x"70"),
  1610 => (x"78",x"c0",x"48",x"d2"),
  1611 => (x"48",x"ce",x"e5",x"c1"),
  1612 => (x"e6",x"c2",x"78",x"c0"),
  1613 => (x"cf",x"fa",x"49",x"ca"),
  1614 => (x"c0",x"4a",x"70",x"87"),
  1615 => (x"fd",x"03",x"aa",x"b7"),
  1616 => (x"48",x"c0",x"87",x"dd"),
  1617 => (x"4d",x"26",x"87",x"c2"),
  1618 => (x"4b",x"26",x"4c",x"26"),
  1619 => (x"00",x"00",x"4f",x"26"),
  1620 => (x"00",x"00",x"00",x"00"),
  1621 => (x"71",x"1e",x"00",x"00"),
  1622 => (x"eb",x"fc",x"49",x"4a"),
  1623 => (x"1e",x"4f",x"26",x"87"),
  1624 => (x"49",x"72",x"4a",x"c0"),
  1625 => (x"e6",x"c1",x"91",x"c4"),
  1626 => (x"79",x"c0",x"81",x"ee"),
  1627 => (x"b7",x"d0",x"82",x"c1"),
  1628 => (x"87",x"ee",x"04",x"aa"),
  1629 => (x"5e",x"0e",x"4f",x"26"),
  1630 => (x"0e",x"5d",x"5c",x"5b"),
  1631 => (x"f7",x"f8",x"4d",x"71"),
  1632 => (x"c4",x"4a",x"75",x"87"),
  1633 => (x"c1",x"92",x"2a",x"b7"),
  1634 => (x"75",x"82",x"ee",x"e6"),
  1635 => (x"c2",x"9c",x"cf",x"4c"),
  1636 => (x"4b",x"49",x"6a",x"94"),
  1637 => (x"9b",x"c3",x"2b",x"74"),
  1638 => (x"30",x"74",x"48",x"c2"),
  1639 => (x"bc",x"ff",x"4c",x"70"),
  1640 => (x"98",x"71",x"48",x"74"),
  1641 => (x"c7",x"f8",x"7a",x"70"),
  1642 => (x"fe",x"48",x"73",x"87"),
  1643 => (x"00",x"00",x"87",x"d8"),
  1644 => (x"00",x"00",x"00",x"00"),
  1645 => (x"00",x"00",x"00",x"00"),
  1646 => (x"00",x"00",x"00",x"00"),
  1647 => (x"00",x"00",x"00",x"00"),
  1648 => (x"00",x"00",x"00",x"00"),
  1649 => (x"00",x"00",x"00",x"00"),
  1650 => (x"00",x"00",x"00",x"00"),
  1651 => (x"00",x"00",x"00",x"00"),
  1652 => (x"00",x"00",x"00",x"00"),
  1653 => (x"00",x"00",x"00",x"00"),
  1654 => (x"00",x"00",x"00",x"00"),
  1655 => (x"00",x"00",x"00",x"00"),
  1656 => (x"00",x"00",x"00",x"00"),
  1657 => (x"00",x"00",x"00",x"00"),
  1658 => (x"00",x"00",x"00",x"00"),
  1659 => (x"ff",x"1e",x"00",x"00"),
  1660 => (x"e1",x"c8",x"48",x"d0"),
  1661 => (x"ff",x"48",x"71",x"78"),
  1662 => (x"c4",x"78",x"08",x"d4"),
  1663 => (x"d4",x"ff",x"48",x"66"),
  1664 => (x"4f",x"26",x"78",x"08"),
  1665 => (x"c4",x"4a",x"71",x"1e"),
  1666 => (x"72",x"1e",x"49",x"66"),
  1667 => (x"87",x"de",x"ff",x"49"),
  1668 => (x"c0",x"48",x"d0",x"ff"),
  1669 => (x"26",x"26",x"78",x"e0"),
  1670 => (x"1e",x"73",x"1e",x"4f"),
  1671 => (x"66",x"c8",x"4b",x"71"),
  1672 => (x"4a",x"73",x"1e",x"49"),
  1673 => (x"49",x"a2",x"e0",x"c1"),
  1674 => (x"26",x"87",x"d9",x"ff"),
  1675 => (x"4d",x"26",x"87",x"c4"),
  1676 => (x"4b",x"26",x"4c",x"26"),
  1677 => (x"71",x"1e",x"4f",x"26"),
  1678 => (x"da",x"1e",x"49",x"4a"),
  1679 => (x"87",x"ee",x"fe",x"49"),
  1680 => (x"49",x"bf",x"66",x"c8"),
  1681 => (x"c4",x"48",x"66",x"c8"),
  1682 => (x"58",x"a6",x"cc",x"80"),
  1683 => (x"ff",x"29",x"b7",x"c8"),
  1684 => (x"78",x"71",x"48",x"d4"),
  1685 => (x"49",x"bf",x"66",x"c8"),
  1686 => (x"71",x"29",x"b7",x"c8"),
  1687 => (x"48",x"d0",x"ff",x"78"),
  1688 => (x"26",x"78",x"e0",x"c0"),
  1689 => (x"ff",x"1e",x"4f",x"26"),
  1690 => (x"ff",x"c3",x"4a",x"d4"),
  1691 => (x"48",x"d0",x"ff",x"7a"),
  1692 => (x"de",x"78",x"e1",x"c0"),
  1693 => (x"d4",x"e6",x"c2",x"7a"),
  1694 => (x"48",x"49",x"7a",x"bf"),
  1695 => (x"7a",x"70",x"28",x"c8"),
  1696 => (x"28",x"d0",x"48",x"71"),
  1697 => (x"48",x"71",x"7a",x"70"),
  1698 => (x"7a",x"70",x"28",x"d8"),
  1699 => (x"c0",x"48",x"d0",x"ff"),
  1700 => (x"4f",x"26",x"78",x"e0"),
  1701 => (x"5c",x"5b",x"5e",x"0e"),
  1702 => (x"4c",x"71",x"0e",x"5d"),
  1703 => (x"bf",x"d4",x"e6",x"c2"),
  1704 => (x"2b",x"74",x"4b",x"4d"),
  1705 => (x"c1",x"9b",x"66",x"d0"),
  1706 => (x"ab",x"66",x"d4",x"83"),
  1707 => (x"c0",x"87",x"c2",x"04"),
  1708 => (x"d0",x"4a",x"74",x"4b"),
  1709 => (x"31",x"72",x"49",x"66"),
  1710 => (x"99",x"75",x"b9",x"ff"),
  1711 => (x"30",x"72",x"48",x"73"),
  1712 => (x"71",x"48",x"4a",x"70"),
  1713 => (x"d8",x"e6",x"c2",x"b0"),
  1714 => (x"87",x"da",x"fe",x"58"),
  1715 => (x"4c",x"26",x"4d",x"26"),
  1716 => (x"4f",x"26",x"4b",x"26"),
  1717 => (x"48",x"d0",x"ff",x"1e"),
  1718 => (x"71",x"78",x"c9",x"c8"),
  1719 => (x"08",x"d4",x"ff",x"48"),
  1720 => (x"1e",x"4f",x"26",x"78"),
  1721 => (x"eb",x"49",x"4a",x"71"),
  1722 => (x"48",x"d0",x"ff",x"87"),
  1723 => (x"4f",x"26",x"78",x"c8"),
  1724 => (x"71",x"1e",x"73",x"1e"),
  1725 => (x"e4",x"e6",x"c2",x"4b"),
  1726 => (x"87",x"c3",x"02",x"bf"),
  1727 => (x"ff",x"87",x"eb",x"c2"),
  1728 => (x"c9",x"c8",x"48",x"d0"),
  1729 => (x"c0",x"49",x"73",x"78"),
  1730 => (x"d4",x"ff",x"b1",x"e0"),
  1731 => (x"c2",x"78",x"71",x"48"),
  1732 => (x"c0",x"48",x"d8",x"e6"),
  1733 => (x"02",x"66",x"c8",x"78"),
  1734 => (x"ff",x"c3",x"87",x"c5"),
  1735 => (x"c0",x"87",x"c2",x"49"),
  1736 => (x"e0",x"e6",x"c2",x"49"),
  1737 => (x"02",x"66",x"cc",x"59"),
  1738 => (x"d5",x"c5",x"87",x"c6"),
  1739 => (x"87",x"c4",x"4a",x"d5"),
  1740 => (x"4a",x"ff",x"ff",x"cf"),
  1741 => (x"5a",x"e4",x"e6",x"c2"),
  1742 => (x"48",x"e4",x"e6",x"c2"),
  1743 => (x"87",x"c4",x"78",x"c1"),
  1744 => (x"4c",x"26",x"4d",x"26"),
  1745 => (x"4f",x"26",x"4b",x"26"),
  1746 => (x"5c",x"5b",x"5e",x"0e"),
  1747 => (x"4a",x"71",x"0e",x"5d"),
  1748 => (x"bf",x"e0",x"e6",x"c2"),
  1749 => (x"02",x"9a",x"72",x"4c"),
  1750 => (x"c8",x"49",x"87",x"cb"),
  1751 => (x"e6",x"eb",x"c1",x"91"),
  1752 => (x"c4",x"83",x"71",x"4b"),
  1753 => (x"e6",x"ef",x"c1",x"87"),
  1754 => (x"13",x"4d",x"c0",x"4b"),
  1755 => (x"c2",x"99",x"74",x"49"),
  1756 => (x"b9",x"bf",x"dc",x"e6"),
  1757 => (x"71",x"48",x"d4",x"ff"),
  1758 => (x"2c",x"b7",x"c1",x"78"),
  1759 => (x"ad",x"b7",x"c8",x"85"),
  1760 => (x"c2",x"87",x"e8",x"04"),
  1761 => (x"48",x"bf",x"d8",x"e6"),
  1762 => (x"e6",x"c2",x"80",x"c8"),
  1763 => (x"ef",x"fe",x"58",x"dc"),
  1764 => (x"1e",x"73",x"1e",x"87"),
  1765 => (x"4a",x"13",x"4b",x"71"),
  1766 => (x"87",x"cb",x"02",x"9a"),
  1767 => (x"e7",x"fe",x"49",x"72"),
  1768 => (x"9a",x"4a",x"13",x"87"),
  1769 => (x"fe",x"87",x"f5",x"05"),
  1770 => (x"c2",x"1e",x"87",x"da"),
  1771 => (x"49",x"bf",x"d8",x"e6"),
  1772 => (x"48",x"d8",x"e6",x"c2"),
  1773 => (x"c4",x"78",x"a1",x"c1"),
  1774 => (x"03",x"a9",x"b7",x"c0"),
  1775 => (x"d4",x"ff",x"87",x"db"),
  1776 => (x"dc",x"e6",x"c2",x"48"),
  1777 => (x"e6",x"c2",x"78",x"bf"),
  1778 => (x"c2",x"49",x"bf",x"d8"),
  1779 => (x"c1",x"48",x"d8",x"e6"),
  1780 => (x"c0",x"c4",x"78",x"a1"),
  1781 => (x"e5",x"04",x"a9",x"b7"),
  1782 => (x"48",x"d0",x"ff",x"87"),
  1783 => (x"e6",x"c2",x"78",x"c8"),
  1784 => (x"78",x"c0",x"48",x"e4"),
  1785 => (x"00",x"00",x"4f",x"26"),
  1786 => (x"00",x"00",x"00",x"00"),
  1787 => (x"00",x"00",x"00",x"00"),
  1788 => (x"00",x"5f",x"5f",x"00"),
  1789 => (x"03",x"00",x"00",x"00"),
  1790 => (x"03",x"03",x"00",x"03"),
  1791 => (x"7f",x"14",x"00",x"00"),
  1792 => (x"7f",x"7f",x"14",x"7f"),
  1793 => (x"24",x"00",x"00",x"14"),
  1794 => (x"3a",x"6b",x"6b",x"2e"),
  1795 => (x"6a",x"4c",x"00",x"12"),
  1796 => (x"56",x"6c",x"18",x"36"),
  1797 => (x"7e",x"30",x"00",x"32"),
  1798 => (x"3a",x"77",x"59",x"4f"),
  1799 => (x"00",x"00",x"40",x"68"),
  1800 => (x"00",x"03",x"07",x"04"),
  1801 => (x"00",x"00",x"00",x"00"),
  1802 => (x"41",x"63",x"3e",x"1c"),
  1803 => (x"00",x"00",x"00",x"00"),
  1804 => (x"1c",x"3e",x"63",x"41"),
  1805 => (x"2a",x"08",x"00",x"00"),
  1806 => (x"3e",x"1c",x"1c",x"3e"),
  1807 => (x"08",x"00",x"08",x"2a"),
  1808 => (x"08",x"3e",x"3e",x"08"),
  1809 => (x"00",x"00",x"00",x"08"),
  1810 => (x"00",x"60",x"e0",x"80"),
  1811 => (x"08",x"00",x"00",x"00"),
  1812 => (x"08",x"08",x"08",x"08"),
  1813 => (x"00",x"00",x"00",x"08"),
  1814 => (x"00",x"60",x"60",x"00"),
  1815 => (x"60",x"40",x"00",x"00"),
  1816 => (x"06",x"0c",x"18",x"30"),
  1817 => (x"3e",x"00",x"01",x"03"),
  1818 => (x"7f",x"4d",x"59",x"7f"),
  1819 => (x"04",x"00",x"00",x"3e"),
  1820 => (x"00",x"7f",x"7f",x"06"),
  1821 => (x"42",x"00",x"00",x"00"),
  1822 => (x"4f",x"59",x"71",x"63"),
  1823 => (x"22",x"00",x"00",x"46"),
  1824 => (x"7f",x"49",x"49",x"63"),
  1825 => (x"1c",x"18",x"00",x"36"),
  1826 => (x"7f",x"7f",x"13",x"16"),
  1827 => (x"27",x"00",x"00",x"10"),
  1828 => (x"7d",x"45",x"45",x"67"),
  1829 => (x"3c",x"00",x"00",x"39"),
  1830 => (x"79",x"49",x"4b",x"7e"),
  1831 => (x"01",x"00",x"00",x"30"),
  1832 => (x"0f",x"79",x"71",x"01"),
  1833 => (x"36",x"00",x"00",x"07"),
  1834 => (x"7f",x"49",x"49",x"7f"),
  1835 => (x"06",x"00",x"00",x"36"),
  1836 => (x"3f",x"69",x"49",x"4f"),
  1837 => (x"00",x"00",x"00",x"1e"),
  1838 => (x"00",x"66",x"66",x"00"),
  1839 => (x"00",x"00",x"00",x"00"),
  1840 => (x"00",x"66",x"e6",x"80"),
  1841 => (x"08",x"00",x"00",x"00"),
  1842 => (x"22",x"14",x"14",x"08"),
  1843 => (x"14",x"00",x"00",x"22"),
  1844 => (x"14",x"14",x"14",x"14"),
  1845 => (x"22",x"00",x"00",x"14"),
  1846 => (x"08",x"14",x"14",x"22"),
  1847 => (x"02",x"00",x"00",x"08"),
  1848 => (x"0f",x"59",x"51",x"03"),
  1849 => (x"7f",x"3e",x"00",x"06"),
  1850 => (x"1f",x"55",x"5d",x"41"),
  1851 => (x"7e",x"00",x"00",x"1e"),
  1852 => (x"7f",x"09",x"09",x"7f"),
  1853 => (x"7f",x"00",x"00",x"7e"),
  1854 => (x"7f",x"49",x"49",x"7f"),
  1855 => (x"1c",x"00",x"00",x"36"),
  1856 => (x"41",x"41",x"63",x"3e"),
  1857 => (x"7f",x"00",x"00",x"41"),
  1858 => (x"3e",x"63",x"41",x"7f"),
  1859 => (x"7f",x"00",x"00",x"1c"),
  1860 => (x"41",x"49",x"49",x"7f"),
  1861 => (x"7f",x"00",x"00",x"41"),
  1862 => (x"01",x"09",x"09",x"7f"),
  1863 => (x"3e",x"00",x"00",x"01"),
  1864 => (x"7b",x"49",x"41",x"7f"),
  1865 => (x"7f",x"00",x"00",x"7a"),
  1866 => (x"7f",x"08",x"08",x"7f"),
  1867 => (x"00",x"00",x"00",x"7f"),
  1868 => (x"41",x"7f",x"7f",x"41"),
  1869 => (x"20",x"00",x"00",x"00"),
  1870 => (x"7f",x"40",x"40",x"60"),
  1871 => (x"7f",x"7f",x"00",x"3f"),
  1872 => (x"63",x"36",x"1c",x"08"),
  1873 => (x"7f",x"00",x"00",x"41"),
  1874 => (x"40",x"40",x"40",x"7f"),
  1875 => (x"7f",x"7f",x"00",x"40"),
  1876 => (x"7f",x"06",x"0c",x"06"),
  1877 => (x"7f",x"7f",x"00",x"7f"),
  1878 => (x"7f",x"18",x"0c",x"06"),
  1879 => (x"3e",x"00",x"00",x"7f"),
  1880 => (x"7f",x"41",x"41",x"7f"),
  1881 => (x"7f",x"00",x"00",x"3e"),
  1882 => (x"0f",x"09",x"09",x"7f"),
  1883 => (x"7f",x"3e",x"00",x"06"),
  1884 => (x"7e",x"7f",x"61",x"41"),
  1885 => (x"7f",x"00",x"00",x"40"),
  1886 => (x"7f",x"19",x"09",x"7f"),
  1887 => (x"26",x"00",x"00",x"66"),
  1888 => (x"7b",x"59",x"4d",x"6f"),
  1889 => (x"01",x"00",x"00",x"32"),
  1890 => (x"01",x"7f",x"7f",x"01"),
  1891 => (x"3f",x"00",x"00",x"01"),
  1892 => (x"7f",x"40",x"40",x"7f"),
  1893 => (x"0f",x"00",x"00",x"3f"),
  1894 => (x"3f",x"70",x"70",x"3f"),
  1895 => (x"7f",x"7f",x"00",x"0f"),
  1896 => (x"7f",x"30",x"18",x"30"),
  1897 => (x"63",x"41",x"00",x"7f"),
  1898 => (x"36",x"1c",x"1c",x"36"),
  1899 => (x"03",x"01",x"41",x"63"),
  1900 => (x"06",x"7c",x"7c",x"06"),
  1901 => (x"71",x"61",x"01",x"03"),
  1902 => (x"43",x"47",x"4d",x"59"),
  1903 => (x"00",x"00",x"00",x"41"),
  1904 => (x"41",x"41",x"7f",x"7f"),
  1905 => (x"03",x"01",x"00",x"00"),
  1906 => (x"30",x"18",x"0c",x"06"),
  1907 => (x"00",x"00",x"40",x"60"),
  1908 => (x"7f",x"7f",x"41",x"41"),
  1909 => (x"0c",x"08",x"00",x"00"),
  1910 => (x"0c",x"06",x"03",x"06"),
  1911 => (x"80",x"80",x"00",x"08"),
  1912 => (x"80",x"80",x"80",x"80"),
  1913 => (x"00",x"00",x"00",x"80"),
  1914 => (x"04",x"07",x"03",x"00"),
  1915 => (x"20",x"00",x"00",x"00"),
  1916 => (x"7c",x"54",x"54",x"74"),
  1917 => (x"7f",x"00",x"00",x"78"),
  1918 => (x"7c",x"44",x"44",x"7f"),
  1919 => (x"38",x"00",x"00",x"38"),
  1920 => (x"44",x"44",x"44",x"7c"),
  1921 => (x"38",x"00",x"00",x"00"),
  1922 => (x"7f",x"44",x"44",x"7c"),
  1923 => (x"38",x"00",x"00",x"7f"),
  1924 => (x"5c",x"54",x"54",x"7c"),
  1925 => (x"04",x"00",x"00",x"18"),
  1926 => (x"05",x"05",x"7f",x"7e"),
  1927 => (x"18",x"00",x"00",x"00"),
  1928 => (x"fc",x"a4",x"a4",x"bc"),
  1929 => (x"7f",x"00",x"00",x"7c"),
  1930 => (x"7c",x"04",x"04",x"7f"),
  1931 => (x"00",x"00",x"00",x"78"),
  1932 => (x"40",x"7d",x"3d",x"00"),
  1933 => (x"80",x"00",x"00",x"00"),
  1934 => (x"7d",x"fd",x"80",x"80"),
  1935 => (x"7f",x"00",x"00",x"00"),
  1936 => (x"6c",x"38",x"10",x"7f"),
  1937 => (x"00",x"00",x"00",x"44"),
  1938 => (x"40",x"7f",x"3f",x"00"),
  1939 => (x"7c",x"7c",x"00",x"00"),
  1940 => (x"7c",x"0c",x"18",x"0c"),
  1941 => (x"7c",x"00",x"00",x"78"),
  1942 => (x"7c",x"04",x"04",x"7c"),
  1943 => (x"38",x"00",x"00",x"78"),
  1944 => (x"7c",x"44",x"44",x"7c"),
  1945 => (x"fc",x"00",x"00",x"38"),
  1946 => (x"3c",x"24",x"24",x"fc"),
  1947 => (x"18",x"00",x"00",x"18"),
  1948 => (x"fc",x"24",x"24",x"3c"),
  1949 => (x"7c",x"00",x"00",x"fc"),
  1950 => (x"0c",x"04",x"04",x"7c"),
  1951 => (x"48",x"00",x"00",x"08"),
  1952 => (x"74",x"54",x"54",x"5c"),
  1953 => (x"04",x"00",x"00",x"20"),
  1954 => (x"44",x"44",x"7f",x"3f"),
  1955 => (x"3c",x"00",x"00",x"00"),
  1956 => (x"7c",x"40",x"40",x"7c"),
  1957 => (x"1c",x"00",x"00",x"7c"),
  1958 => (x"3c",x"60",x"60",x"3c"),
  1959 => (x"7c",x"3c",x"00",x"1c"),
  1960 => (x"7c",x"60",x"30",x"60"),
  1961 => (x"6c",x"44",x"00",x"3c"),
  1962 => (x"6c",x"38",x"10",x"38"),
  1963 => (x"1c",x"00",x"00",x"44"),
  1964 => (x"3c",x"60",x"e0",x"bc"),
  1965 => (x"44",x"00",x"00",x"1c"),
  1966 => (x"4c",x"5c",x"74",x"64"),
  1967 => (x"08",x"00",x"00",x"44"),
  1968 => (x"41",x"77",x"3e",x"08"),
  1969 => (x"00",x"00",x"00",x"41"),
  1970 => (x"00",x"7f",x"7f",x"00"),
  1971 => (x"41",x"00",x"00",x"00"),
  1972 => (x"08",x"3e",x"77",x"41"),
  1973 => (x"01",x"02",x"00",x"08"),
  1974 => (x"02",x"02",x"03",x"01"),
  1975 => (x"7f",x"7f",x"00",x"01"),
  1976 => (x"7f",x"7f",x"7f",x"7f"),
  1977 => (x"08",x"08",x"00",x"7f"),
  1978 => (x"3e",x"3e",x"1c",x"1c"),
  1979 => (x"7f",x"7f",x"7f",x"7f"),
  1980 => (x"1c",x"1c",x"3e",x"3e"),
  1981 => (x"10",x"00",x"08",x"08"),
  1982 => (x"18",x"7c",x"7c",x"18"),
  1983 => (x"10",x"00",x"00",x"10"),
  1984 => (x"30",x"7c",x"7c",x"30"),
  1985 => (x"30",x"10",x"00",x"10"),
  1986 => (x"1e",x"78",x"60",x"60"),
  1987 => (x"66",x"42",x"00",x"06"),
  1988 => (x"66",x"3c",x"18",x"3c"),
  1989 => (x"38",x"78",x"00",x"42"),
  1990 => (x"6c",x"c6",x"c2",x"6a"),
  1991 => (x"00",x"60",x"00",x"38"),
  1992 => (x"00",x"00",x"60",x"00"),
  1993 => (x"5e",x"0e",x"00",x"60"),
  1994 => (x"0e",x"5d",x"5c",x"5b"),
  1995 => (x"c2",x"4c",x"71",x"1e"),
  1996 => (x"4d",x"bf",x"f5",x"e6"),
  1997 => (x"1e",x"c0",x"4b",x"c0"),
  1998 => (x"c7",x"02",x"ab",x"74"),
  1999 => (x"48",x"a6",x"c4",x"87"),
  2000 => (x"87",x"c5",x"78",x"c0"),
  2001 => (x"c1",x"48",x"a6",x"c4"),
  2002 => (x"1e",x"66",x"c4",x"78"),
  2003 => (x"df",x"ee",x"49",x"73"),
  2004 => (x"c0",x"86",x"c8",x"87"),
  2005 => (x"ef",x"ef",x"49",x"e0"),
  2006 => (x"4a",x"a5",x"c4",x"87"),
  2007 => (x"f0",x"f0",x"49",x"6a"),
  2008 => (x"87",x"c6",x"f1",x"87"),
  2009 => (x"83",x"c1",x"85",x"cb"),
  2010 => (x"04",x"ab",x"b7",x"c8"),
  2011 => (x"26",x"87",x"c7",x"ff"),
  2012 => (x"4c",x"26",x"4d",x"26"),
  2013 => (x"4f",x"26",x"4b",x"26"),
  2014 => (x"c2",x"4a",x"71",x"1e"),
  2015 => (x"c2",x"5a",x"f9",x"e6"),
  2016 => (x"c7",x"48",x"f9",x"e6"),
  2017 => (x"dd",x"fe",x"49",x"78"),
  2018 => (x"1e",x"4f",x"26",x"87"),
  2019 => (x"4a",x"71",x"1e",x"73"),
  2020 => (x"03",x"aa",x"b7",x"c0"),
  2021 => (x"cd",x"c2",x"87",x"d3"),
  2022 => (x"c4",x"05",x"bf",x"d8"),
  2023 => (x"c2",x"4b",x"c1",x"87"),
  2024 => (x"c2",x"4b",x"c0",x"87"),
  2025 => (x"c4",x"5b",x"dc",x"cd"),
  2026 => (x"dc",x"cd",x"c2",x"87"),
  2027 => (x"d8",x"cd",x"c2",x"5a"),
  2028 => (x"9a",x"c1",x"4a",x"bf"),
  2029 => (x"49",x"a2",x"c0",x"c1"),
  2030 => (x"fc",x"87",x"e8",x"ec"),
  2031 => (x"d8",x"cd",x"c2",x"48"),
  2032 => (x"ef",x"fe",x"78",x"bf"),
  2033 => (x"5b",x"5e",x"0e",x"87"),
  2034 => (x"71",x"0e",x"5d",x"5c"),
  2035 => (x"f8",x"4a",x"6b",x"4b"),
  2036 => (x"c7",x"4d",x"c0",x"c4"),
  2037 => (x"d0",x"4c",x"c0",x"fc"),
  2038 => (x"99",x"c2",x"49",x"66"),
  2039 => (x"d4",x"87",x"cf",x"02"),
  2040 => (x"09",x"c0",x"49",x"66"),
  2041 => (x"c8",x"4c",x"71",x"89"),
  2042 => (x"8a",x"66",x"d4",x"34"),
  2043 => (x"66",x"d0",x"87",x"d7"),
  2044 => (x"02",x"99",x"c1",x"49"),
  2045 => (x"66",x"d4",x"87",x"ca"),
  2046 => (x"d4",x"35",x"c8",x"4d"),
  2047 => (x"87",x"c5",x"82",x"66"),
  2048 => (x"b7",x"c4",x"92",x"cf"),
  2049 => (x"aa",x"b7",x"75",x"2a"),
  2050 => (x"4a",x"87",x"c1",x"03"),
  2051 => (x"06",x"aa",x"b7",x"74"),
  2052 => (x"72",x"4a",x"87",x"c1"),
  2053 => (x"87",x"d8",x"fd",x"7b"),
  2054 => (x"d8",x"cd",x"c2",x"1e"),
  2055 => (x"f5",x"e4",x"49",x"bf"),
  2056 => (x"ed",x"e6",x"c2",x"87"),
  2057 => (x"78",x"bf",x"e8",x"48"),
  2058 => (x"48",x"e9",x"e6",x"c2"),
  2059 => (x"c2",x"78",x"bf",x"ec"),
  2060 => (x"4a",x"bf",x"ed",x"e6"),
  2061 => (x"99",x"ff",x"c3",x"49"),
  2062 => (x"72",x"2a",x"b7",x"c8"),
  2063 => (x"c2",x"b0",x"71",x"48"),
  2064 => (x"26",x"58",x"f5",x"e6"),
  2065 => (x"5b",x"5e",x"0e",x"4f"),
  2066 => (x"71",x"0e",x"5d",x"5c"),
  2067 => (x"87",x"c8",x"ff",x"4b"),
  2068 => (x"48",x"e8",x"e6",x"c2"),
  2069 => (x"49",x"73",x"50",x"c0"),
  2070 => (x"70",x"87",x"db",x"e4"),
  2071 => (x"9c",x"c2",x"4c",x"49"),
  2072 => (x"cb",x"49",x"ee",x"cb"),
  2073 => (x"49",x"70",x"87",x"fa"),
  2074 => (x"e8",x"e6",x"c2",x"4d"),
  2075 => (x"c1",x"05",x"bf",x"97"),
  2076 => (x"66",x"d0",x"87",x"e2"),
  2077 => (x"f1",x"e6",x"c2",x"49"),
  2078 => (x"d6",x"05",x"99",x"bf"),
  2079 => (x"49",x"66",x"d4",x"87"),
  2080 => (x"bf",x"e9",x"e6",x"c2"),
  2081 => (x"87",x"cb",x"05",x"99"),
  2082 => (x"e9",x"e3",x"49",x"73"),
  2083 => (x"02",x"98",x"70",x"87"),
  2084 => (x"c1",x"87",x"c1",x"c1"),
  2085 => (x"87",x"c0",x"fe",x"4c"),
  2086 => (x"cf",x"cb",x"49",x"75"),
  2087 => (x"02",x"98",x"70",x"87"),
  2088 => (x"e6",x"c2",x"87",x"c6"),
  2089 => (x"50",x"c1",x"48",x"e8"),
  2090 => (x"97",x"e8",x"e6",x"c2"),
  2091 => (x"e3",x"c0",x"05",x"bf"),
  2092 => (x"f1",x"e6",x"c2",x"87"),
  2093 => (x"66",x"d0",x"49",x"bf"),
  2094 => (x"d6",x"ff",x"05",x"99"),
  2095 => (x"e9",x"e6",x"c2",x"87"),
  2096 => (x"66",x"d4",x"49",x"bf"),
  2097 => (x"ca",x"ff",x"05",x"99"),
  2098 => (x"e2",x"49",x"73",x"87"),
  2099 => (x"98",x"70",x"87",x"e8"),
  2100 => (x"87",x"ff",x"fe",x"05"),
  2101 => (x"d7",x"fa",x"48",x"74"),
  2102 => (x"5b",x"5e",x"0e",x"87"),
  2103 => (x"f4",x"0e",x"5d",x"5c"),
  2104 => (x"4c",x"4d",x"c0",x"86"),
  2105 => (x"c4",x"7e",x"bf",x"ec"),
  2106 => (x"e6",x"c2",x"48",x"a6"),
  2107 => (x"c1",x"78",x"bf",x"f5"),
  2108 => (x"c7",x"1e",x"c0",x"1e"),
  2109 => (x"87",x"cd",x"fd",x"49"),
  2110 => (x"98",x"70",x"86",x"c8"),
  2111 => (x"ff",x"87",x"cd",x"02"),
  2112 => (x"87",x"c7",x"fa",x"49"),
  2113 => (x"e1",x"49",x"da",x"c1"),
  2114 => (x"4d",x"c1",x"87",x"ec"),
  2115 => (x"97",x"e8",x"e6",x"c2"),
  2116 => (x"87",x"c3",x"02",x"bf"),
  2117 => (x"c2",x"87",x"ee",x"c9"),
  2118 => (x"4b",x"bf",x"ed",x"e6"),
  2119 => (x"bf",x"d8",x"cd",x"c2"),
  2120 => (x"87",x"d9",x"c1",x"05"),
  2121 => (x"c8",x"48",x"a6",x"c4"),
  2122 => (x"c2",x"78",x"c0",x"c0"),
  2123 => (x"6e",x"7e",x"dd",x"d4"),
  2124 => (x"6e",x"49",x"bf",x"97"),
  2125 => (x"70",x"80",x"c1",x"48"),
  2126 => (x"f9",x"e0",x"71",x"7e"),
  2127 => (x"02",x"98",x"70",x"87"),
  2128 => (x"66",x"c4",x"87",x"c3"),
  2129 => (x"48",x"66",x"c4",x"b3"),
  2130 => (x"c8",x"28",x"b7",x"c1"),
  2131 => (x"98",x"70",x"58",x"a6"),
  2132 => (x"87",x"db",x"ff",x"05"),
  2133 => (x"e0",x"49",x"fd",x"c3"),
  2134 => (x"fa",x"c3",x"87",x"dc"),
  2135 => (x"87",x"d6",x"e0",x"49"),
  2136 => (x"ff",x"c3",x"49",x"73"),
  2137 => (x"c0",x"1e",x"71",x"99"),
  2138 => (x"87",x"c6",x"c9",x"49"),
  2139 => (x"b7",x"c8",x"49",x"73"),
  2140 => (x"c1",x"1e",x"71",x"29"),
  2141 => (x"87",x"fa",x"c8",x"49"),
  2142 => (x"c1",x"c6",x"86",x"c8"),
  2143 => (x"f1",x"e6",x"c2",x"87"),
  2144 => (x"02",x"9b",x"4b",x"bf"),
  2145 => (x"cd",x"c2",x"87",x"dd"),
  2146 => (x"c7",x"49",x"bf",x"d4"),
  2147 => (x"98",x"70",x"87",x"de"),
  2148 => (x"c0",x"87",x"c4",x"05"),
  2149 => (x"c2",x"87",x"d2",x"4b"),
  2150 => (x"c3",x"c7",x"49",x"e0"),
  2151 => (x"d8",x"cd",x"c2",x"87"),
  2152 => (x"c2",x"87",x"c6",x"58"),
  2153 => (x"c0",x"48",x"d4",x"cd"),
  2154 => (x"c2",x"49",x"73",x"78"),
  2155 => (x"87",x"ce",x"05",x"99"),
  2156 => (x"ff",x"49",x"eb",x"c3"),
  2157 => (x"70",x"87",x"ff",x"de"),
  2158 => (x"02",x"99",x"c2",x"49"),
  2159 => (x"4c",x"fb",x"87",x"c2"),
  2160 => (x"99",x"c1",x"49",x"73"),
  2161 => (x"c3",x"87",x"ce",x"05"),
  2162 => (x"de",x"ff",x"49",x"f4"),
  2163 => (x"49",x"70",x"87",x"e8"),
  2164 => (x"c2",x"02",x"99",x"c2"),
  2165 => (x"73",x"4c",x"fa",x"87"),
  2166 => (x"05",x"99",x"c8",x"49"),
  2167 => (x"f5",x"c3",x"87",x"ce"),
  2168 => (x"d1",x"de",x"ff",x"49"),
  2169 => (x"c2",x"49",x"70",x"87"),
  2170 => (x"87",x"d5",x"02",x"99"),
  2171 => (x"bf",x"f9",x"e6",x"c2"),
  2172 => (x"48",x"87",x"ca",x"02"),
  2173 => (x"e6",x"c2",x"88",x"c1"),
  2174 => (x"c2",x"c0",x"58",x"fd"),
  2175 => (x"c1",x"4c",x"ff",x"87"),
  2176 => (x"c4",x"49",x"73",x"4d"),
  2177 => (x"87",x"ce",x"05",x"99"),
  2178 => (x"ff",x"49",x"f2",x"c3"),
  2179 => (x"70",x"87",x"e7",x"dd"),
  2180 => (x"02",x"99",x"c2",x"49"),
  2181 => (x"e6",x"c2",x"87",x"dc"),
  2182 => (x"48",x"7e",x"bf",x"f9"),
  2183 => (x"03",x"a8",x"b7",x"c7"),
  2184 => (x"6e",x"87",x"cb",x"c0"),
  2185 => (x"c2",x"80",x"c1",x"48"),
  2186 => (x"c0",x"58",x"fd",x"e6"),
  2187 => (x"4c",x"fe",x"87",x"c2"),
  2188 => (x"fd",x"c3",x"4d",x"c1"),
  2189 => (x"fd",x"dc",x"ff",x"49"),
  2190 => (x"c2",x"49",x"70",x"87"),
  2191 => (x"d5",x"c0",x"02",x"99"),
  2192 => (x"f9",x"e6",x"c2",x"87"),
  2193 => (x"c9",x"c0",x"02",x"bf"),
  2194 => (x"f9",x"e6",x"c2",x"87"),
  2195 => (x"c0",x"78",x"c0",x"48"),
  2196 => (x"4c",x"fd",x"87",x"c2"),
  2197 => (x"fa",x"c3",x"4d",x"c1"),
  2198 => (x"d9",x"dc",x"ff",x"49"),
  2199 => (x"c2",x"49",x"70",x"87"),
  2200 => (x"d9",x"c0",x"02",x"99"),
  2201 => (x"f9",x"e6",x"c2",x"87"),
  2202 => (x"b7",x"c7",x"48",x"bf"),
  2203 => (x"c9",x"c0",x"03",x"a8"),
  2204 => (x"f9",x"e6",x"c2",x"87"),
  2205 => (x"c0",x"78",x"c7",x"48"),
  2206 => (x"4c",x"fc",x"87",x"c2"),
  2207 => (x"b7",x"c0",x"4d",x"c1"),
  2208 => (x"d1",x"c0",x"03",x"ac"),
  2209 => (x"4a",x"66",x"c4",x"87"),
  2210 => (x"6a",x"82",x"d8",x"c1"),
  2211 => (x"87",x"c6",x"c0",x"02"),
  2212 => (x"49",x"74",x"4b",x"6a"),
  2213 => (x"1e",x"c0",x"0f",x"73"),
  2214 => (x"c1",x"1e",x"f0",x"c3"),
  2215 => (x"e4",x"f6",x"49",x"da"),
  2216 => (x"70",x"86",x"c8",x"87"),
  2217 => (x"e2",x"c0",x"02",x"98"),
  2218 => (x"48",x"a6",x"c8",x"87"),
  2219 => (x"bf",x"f9",x"e6",x"c2"),
  2220 => (x"49",x"66",x"c8",x"78"),
  2221 => (x"66",x"c4",x"91",x"cb"),
  2222 => (x"70",x"80",x"71",x"48"),
  2223 => (x"02",x"bf",x"6e",x"7e"),
  2224 => (x"6e",x"87",x"c8",x"c0"),
  2225 => (x"66",x"c8",x"4b",x"bf"),
  2226 => (x"75",x"0f",x"73",x"49"),
  2227 => (x"c8",x"c0",x"02",x"9d"),
  2228 => (x"f9",x"e6",x"c2",x"87"),
  2229 => (x"cd",x"f1",x"49",x"bf"),
  2230 => (x"dc",x"cd",x"c2",x"87"),
  2231 => (x"dd",x"c0",x"02",x"bf"),
  2232 => (x"c7",x"c2",x"49",x"87"),
  2233 => (x"02",x"98",x"70",x"87"),
  2234 => (x"c2",x"87",x"d3",x"c0"),
  2235 => (x"49",x"bf",x"f9",x"e6"),
  2236 => (x"c0",x"87",x"f3",x"f0"),
  2237 => (x"87",x"d3",x"f2",x"49"),
  2238 => (x"48",x"dc",x"cd",x"c2"),
  2239 => (x"8e",x"f4",x"78",x"c0"),
  2240 => (x"0e",x"87",x"ed",x"f1"),
  2241 => (x"5d",x"5c",x"5b",x"5e"),
  2242 => (x"4c",x"71",x"1e",x"0e"),
  2243 => (x"bf",x"f5",x"e6",x"c2"),
  2244 => (x"a1",x"cd",x"c1",x"49"),
  2245 => (x"81",x"d1",x"c1",x"4d"),
  2246 => (x"9c",x"74",x"7e",x"69"),
  2247 => (x"c4",x"87",x"cf",x"02"),
  2248 => (x"7b",x"74",x"4b",x"a5"),
  2249 => (x"bf",x"f5",x"e6",x"c2"),
  2250 => (x"87",x"cc",x"f1",x"49"),
  2251 => (x"9c",x"74",x"7b",x"6e"),
  2252 => (x"c0",x"87",x"c4",x"05"),
  2253 => (x"c1",x"87",x"c2",x"4b"),
  2254 => (x"f1",x"49",x"73",x"4b"),
  2255 => (x"66",x"d4",x"87",x"cd"),
  2256 => (x"49",x"87",x"c7",x"02"),
  2257 => (x"4a",x"70",x"87",x"da"),
  2258 => (x"4a",x"c0",x"87",x"c2"),
  2259 => (x"5a",x"e0",x"cd",x"c2"),
  2260 => (x"87",x"dc",x"f0",x"26"),
  2261 => (x"00",x"00",x"00",x"00"),
  2262 => (x"00",x"00",x"00",x"00"),
  2263 => (x"00",x"00",x"00",x"00"),
  2264 => (x"ff",x"4a",x"71",x"1e"),
  2265 => (x"72",x"49",x"bf",x"c8"),
  2266 => (x"4f",x"26",x"48",x"a1"),
  2267 => (x"bf",x"c8",x"ff",x"1e"),
  2268 => (x"c0",x"c0",x"fe",x"89"),
  2269 => (x"a9",x"c0",x"c0",x"c0"),
  2270 => (x"c0",x"87",x"c4",x"01"),
  2271 => (x"c1",x"87",x"c2",x"4a"),
  2272 => (x"26",x"48",x"72",x"4a"),
  2273 => (x"ce",x"c2",x"1e",x"4f"),
  2274 => (x"c1",x"49",x"bf",x"ee"),
  2275 => (x"f2",x"ce",x"c2",x"b9"),
  2276 => (x"48",x"d4",x"ff",x"59"),
  2277 => (x"ff",x"78",x"ff",x"c3"),
  2278 => (x"e1",x"c0",x"48",x"d0"),
  2279 => (x"48",x"d4",x"ff",x"78"),
  2280 => (x"31",x"c4",x"78",x"c1"),
  2281 => (x"d0",x"ff",x"78",x"71"),
  2282 => (x"78",x"e0",x"c0",x"48"),
  2283 => (x"00",x"00",x"4f",x"26"),
  2284 => (x"5e",x"0e",x"00",x"00"),
  2285 => (x"0e",x"5d",x"5c",x"5b"),
  2286 => (x"bf",x"ec",x"4d",x"71"),
  2287 => (x"ff",x"49",x"c5",x"4b"),
  2288 => (x"70",x"87",x"f3",x"d6"),
  2289 => (x"87",x"c7",x"05",x"98"),
  2290 => (x"99",x"c2",x"49",x"73"),
  2291 => (x"c2",x"87",x"c7",x"02"),
  2292 => (x"c2",x"48",x"ed",x"d4"),
  2293 => (x"49",x"c6",x"78",x"c0"),
  2294 => (x"87",x"da",x"d6",x"ff"),
  2295 => (x"c7",x"05",x"98",x"70"),
  2296 => (x"c4",x"49",x"73",x"87"),
  2297 => (x"87",x"c7",x"02",x"99"),
  2298 => (x"48",x"ed",x"d4",x"c2"),
  2299 => (x"c4",x"78",x"f0",x"c0"),
  2300 => (x"c1",x"d6",x"ff",x"49"),
  2301 => (x"05",x"98",x"70",x"87"),
  2302 => (x"49",x"73",x"87",x"c7"),
  2303 => (x"c6",x"02",x"99",x"c8"),
  2304 => (x"ed",x"d4",x"c2",x"87"),
  2305 => (x"cc",x"78",x"cc",x"48"),
  2306 => (x"e9",x"d5",x"ff",x"49"),
  2307 => (x"05",x"98",x"70",x"87"),
  2308 => (x"49",x"73",x"87",x"c7"),
  2309 => (x"c6",x"02",x"99",x"d0"),
  2310 => (x"ed",x"d4",x"c2",x"87"),
  2311 => (x"d0",x"78",x"c8",x"48"),
  2312 => (x"49",x"75",x"1e",x"66"),
  2313 => (x"87",x"f1",x"d7",x"ff"),
  2314 => (x"bf",x"ed",x"d4",x"c2"),
  2315 => (x"1e",x"66",x"d8",x"1e"),
  2316 => (x"93",x"c2",x"4b",x"75"),
  2317 => (x"94",x"c8",x"4c",x"75"),
  2318 => (x"84",x"fd",x"e6",x"c2"),
  2319 => (x"c4",x"ee",x"49",x"6c"),
  2320 => (x"c2",x"7c",x"70",x"87"),
  2321 => (x"1e",x"bf",x"ed",x"d4"),
  2322 => (x"49",x"66",x"e0",x"c0"),
  2323 => (x"71",x"29",x"b7",x"c2"),
  2324 => (x"c2",x"93",x"c4",x"1e"),
  2325 => (x"6b",x"83",x"c1",x"e7"),
  2326 => (x"87",x"e9",x"ed",x"49"),
  2327 => (x"e6",x"c2",x"7b",x"70"),
  2328 => (x"49",x"75",x"1e",x"fd"),
  2329 => (x"87",x"ce",x"d7",x"ff"),
  2330 => (x"4d",x"26",x"8e",x"e8"),
  2331 => (x"4b",x"26",x"4c",x"26"),
  2332 => (x"73",x"1e",x"4f",x"26"),
  2333 => (x"df",x"dc",x"c1",x"1e"),
  2334 => (x"c2",x"50",x"c0",x"48"),
  2335 => (x"c2",x"48",x"f0",x"d4"),
  2336 => (x"c2",x"78",x"c0",x"c0"),
  2337 => (x"48",x"bf",x"d4",x"e6"),
  2338 => (x"e6",x"c2",x"b0",x"c1"),
  2339 => (x"d7",x"ff",x"58",x"d8"),
  2340 => (x"d3",x"c2",x"87",x"d4"),
  2341 => (x"e3",x"fe",x"49",x"ee"),
  2342 => (x"4b",x"70",x"87",x"c2"),
  2343 => (x"bf",x"d4",x"e6",x"c2"),
  2344 => (x"c2",x"98",x"fe",x"48"),
  2345 => (x"ff",x"58",x"d8",x"e6"),
  2346 => (x"73",x"87",x"fb",x"d6"),
  2347 => (x"87",x"c7",x"05",x"9b"),
  2348 => (x"48",x"fa",x"d3",x"c2"),
  2349 => (x"c2",x"87",x"f4",x"c0"),
  2350 => (x"48",x"bf",x"d4",x"e6"),
  2351 => (x"e6",x"c2",x"b0",x"c1"),
  2352 => (x"d6",x"ff",x"58",x"d8"),
  2353 => (x"d4",x"c2",x"87",x"e0"),
  2354 => (x"78",x"c1",x"48",x"f0"),
  2355 => (x"48",x"df",x"dc",x"c1"),
  2356 => (x"d4",x"c2",x"50",x"c1"),
  2357 => (x"e2",x"fe",x"49",x"d1"),
  2358 => (x"e6",x"c2",x"87",x"c2"),
  2359 => (x"fe",x"48",x"bf",x"d4"),
  2360 => (x"d8",x"e6",x"c2",x"98"),
  2361 => (x"fd",x"d5",x"ff",x"58"),
  2362 => (x"fe",x"48",x"c0",x"87"),
  2363 => (x"45",x"56",x"87",x"c0"),
  2364 => (x"45",x"52",x"54",x"43"),
  2365 => (x"49",x"42",x"20",x"58"),
  2366 => (x"45",x"56",x"00",x"4e"),
  2367 => (x"45",x"52",x"54",x"43"),
  2368 => (x"49",x"42",x"2e",x"58"),
  2369 => (x"6f",x"6e",x"20",x"4e"),
  2370 => (x"6f",x"66",x"20",x"74"),
  2371 => (x"21",x"64",x"6e",x"75"),
  2372 => (x"54",x"55",x"41",x"00"),
  2373 => (x"4f",x"4f",x"42",x"4f"),
  2374 => (x"43",x"45",x"56",x"54"),
  2375 => (x"14",x"12",x"58",x"00"),
  2376 => (x"1c",x"1b",x"1d",x"11"),
  2377 => (x"49",x"4a",x"59",x"23"),
  2378 => (x"eb",x"f2",x"f5",x"41"),
  2379 => (x"00",x"00",x"80",x"f4"),
  2380 => (x"00",x"00",x"80",x"00"),
		others => (others => x"00")
	);
	signal q1_local : word_t;

	-- Altera Quartus attributes
	attribute ramstyle: string;
	attribute ramstyle of ram: signal is "no_rw_check";

begin  -- rtl

	addr1 <= to_integer(unsigned(addr(ADDR_WIDTH-1 downto 0)));

	-- Reorganize the read data from the RAM to match the output
	q(7 downto 0) <= q1_local(3);
	q(15 downto 8) <= q1_local(2);
	q(23 downto 16) <= q1_local(1);
	q(31 downto 24) <= q1_local(0);

	process(clk)
	begin
		if(rising_edge(clk)) then 
			if(we = '1') then
				-- edit this code if using other than four bytes per word
				if (bytesel(3) = '1') then
					ram(addr1)(3) <= d(7 downto 0);
				end if;
				if (bytesel(2) = '1') then
					ram(addr1)(2) <= d(15 downto 8);
				end if;
				if (bytesel(1) = '1') then
					ram(addr1)(1) <= d(23 downto 16);
				end if;
				if (bytesel(0) = '1') then
					ram(addr1)(0) <= d(31 downto 24);
				end if;
			end if;
			q1_local <= ram(addr1);
		end if;
	end process;
  
end rtl;

