
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity controller_rom2 is
generic
	(
		ADDR_WIDTH : integer := 15 -- Specify your actual ROM size to save LEs and unnecessary block RAM usage.
	);
port (
	clk : in std_logic;
	reset_n : in std_logic := '1';
	addr : in std_logic_vector(ADDR_WIDTH-1 downto 0);
	q : out std_logic_vector(31 downto 0);
	-- Allow writes - defaults supplied to simplify projects that don't need to write.
	d : in std_logic_vector(31 downto 0) := X"00000000";
	we : in std_logic := '0';
	bytesel : in std_logic_vector(3 downto 0) := "1111"
);
end entity;

architecture rtl of controller_rom2 is

	signal addr1 : integer range 0 to 2**ADDR_WIDTH-1;

	--  build up 2D array to hold the memory
	type word_t is array (0 to 3) of std_logic_vector(7 downto 0);
	type ram_t is array (0 to 2 ** ADDR_WIDTH - 1) of word_t;

	signal ram : ram_t:=
	(

     0 => (x"b7",x"c4",x"92",x"cf"),
     1 => (x"aa",x"b7",x"75",x"2a"),
     2 => (x"4a",x"87",x"c1",x"03"),
     3 => (x"06",x"aa",x"b7",x"74"),
     4 => (x"72",x"4a",x"87",x"c1"),
     5 => (x"87",x"d8",x"fd",x"7b"),
     6 => (x"d8",x"cd",x"c2",x"1e"),
     7 => (x"f5",x"e4",x"49",x"bf"),
     8 => (x"ed",x"e6",x"c2",x"87"),
     9 => (x"78",x"bf",x"e8",x"48"),
    10 => (x"48",x"e9",x"e6",x"c2"),
    11 => (x"c2",x"78",x"bf",x"ec"),
    12 => (x"4a",x"bf",x"ed",x"e6"),
    13 => (x"99",x"ff",x"c3",x"49"),
    14 => (x"72",x"2a",x"b7",x"c8"),
    15 => (x"c2",x"b0",x"71",x"48"),
    16 => (x"26",x"58",x"f5",x"e6"),
    17 => (x"5b",x"5e",x"0e",x"4f"),
    18 => (x"71",x"0e",x"5d",x"5c"),
    19 => (x"87",x"c8",x"ff",x"4b"),
    20 => (x"48",x"e8",x"e6",x"c2"),
    21 => (x"49",x"73",x"50",x"c0"),
    22 => (x"70",x"87",x"db",x"e4"),
    23 => (x"9c",x"c2",x"4c",x"49"),
    24 => (x"cb",x"49",x"ee",x"cb"),
    25 => (x"49",x"70",x"87",x"fa"),
    26 => (x"e8",x"e6",x"c2",x"4d"),
    27 => (x"c1",x"05",x"bf",x"97"),
    28 => (x"66",x"d0",x"87",x"e2"),
    29 => (x"f1",x"e6",x"c2",x"49"),
    30 => (x"d6",x"05",x"99",x"bf"),
    31 => (x"49",x"66",x"d4",x"87"),
    32 => (x"bf",x"e9",x"e6",x"c2"),
    33 => (x"87",x"cb",x"05",x"99"),
    34 => (x"e9",x"e3",x"49",x"73"),
    35 => (x"02",x"98",x"70",x"87"),
    36 => (x"c1",x"87",x"c1",x"c1"),
    37 => (x"87",x"c0",x"fe",x"4c"),
    38 => (x"cf",x"cb",x"49",x"75"),
    39 => (x"02",x"98",x"70",x"87"),
    40 => (x"e6",x"c2",x"87",x"c6"),
    41 => (x"50",x"c1",x"48",x"e8"),
    42 => (x"97",x"e8",x"e6",x"c2"),
    43 => (x"e3",x"c0",x"05",x"bf"),
    44 => (x"f1",x"e6",x"c2",x"87"),
    45 => (x"66",x"d0",x"49",x"bf"),
    46 => (x"d6",x"ff",x"05",x"99"),
    47 => (x"e9",x"e6",x"c2",x"87"),
    48 => (x"66",x"d4",x"49",x"bf"),
    49 => (x"ca",x"ff",x"05",x"99"),
    50 => (x"e2",x"49",x"73",x"87"),
    51 => (x"98",x"70",x"87",x"e8"),
    52 => (x"87",x"ff",x"fe",x"05"),
    53 => (x"d7",x"fa",x"48",x"74"),
    54 => (x"5b",x"5e",x"0e",x"87"),
    55 => (x"f4",x"0e",x"5d",x"5c"),
    56 => (x"4c",x"4d",x"c0",x"86"),
    57 => (x"c4",x"7e",x"bf",x"ec"),
    58 => (x"e6",x"c2",x"48",x"a6"),
    59 => (x"c1",x"78",x"bf",x"f5"),
    60 => (x"c7",x"1e",x"c0",x"1e"),
    61 => (x"87",x"cd",x"fd",x"49"),
    62 => (x"98",x"70",x"86",x"c8"),
    63 => (x"ff",x"87",x"cd",x"02"),
    64 => (x"87",x"c7",x"fa",x"49"),
    65 => (x"e1",x"49",x"da",x"c1"),
    66 => (x"4d",x"c1",x"87",x"ec"),
    67 => (x"97",x"e8",x"e6",x"c2"),
    68 => (x"87",x"c3",x"02",x"bf"),
    69 => (x"c2",x"87",x"ee",x"c9"),
    70 => (x"4b",x"bf",x"ed",x"e6"),
    71 => (x"bf",x"d8",x"cd",x"c2"),
    72 => (x"87",x"d9",x"c1",x"05"),
    73 => (x"c8",x"48",x"a6",x"c4"),
    74 => (x"c2",x"78",x"c0",x"c0"),
    75 => (x"6e",x"7e",x"dd",x"d4"),
    76 => (x"6e",x"49",x"bf",x"97"),
    77 => (x"70",x"80",x"c1",x"48"),
    78 => (x"f9",x"e0",x"71",x"7e"),
    79 => (x"02",x"98",x"70",x"87"),
    80 => (x"66",x"c4",x"87",x"c3"),
    81 => (x"48",x"66",x"c4",x"b3"),
    82 => (x"c8",x"28",x"b7",x"c1"),
    83 => (x"98",x"70",x"58",x"a6"),
    84 => (x"87",x"db",x"ff",x"05"),
    85 => (x"e0",x"49",x"fd",x"c3"),
    86 => (x"fa",x"c3",x"87",x"dc"),
    87 => (x"87",x"d6",x"e0",x"49"),
    88 => (x"ff",x"c3",x"49",x"73"),
    89 => (x"c0",x"1e",x"71",x"99"),
    90 => (x"87",x"c6",x"c9",x"49"),
    91 => (x"b7",x"c8",x"49",x"73"),
    92 => (x"c1",x"1e",x"71",x"29"),
    93 => (x"87",x"fa",x"c8",x"49"),
    94 => (x"c1",x"c6",x"86",x"c8"),
    95 => (x"f1",x"e6",x"c2",x"87"),
    96 => (x"02",x"9b",x"4b",x"bf"),
    97 => (x"cd",x"c2",x"87",x"dd"),
    98 => (x"c7",x"49",x"bf",x"d4"),
    99 => (x"98",x"70",x"87",x"de"),
   100 => (x"c0",x"87",x"c4",x"05"),
   101 => (x"c2",x"87",x"d2",x"4b"),
   102 => (x"c3",x"c7",x"49",x"e0"),
   103 => (x"d8",x"cd",x"c2",x"87"),
   104 => (x"c2",x"87",x"c6",x"58"),
   105 => (x"c0",x"48",x"d4",x"cd"),
   106 => (x"c2",x"49",x"73",x"78"),
   107 => (x"87",x"ce",x"05",x"99"),
   108 => (x"ff",x"49",x"eb",x"c3"),
   109 => (x"70",x"87",x"ff",x"de"),
   110 => (x"02",x"99",x"c2",x"49"),
   111 => (x"4c",x"fb",x"87",x"c2"),
   112 => (x"99",x"c1",x"49",x"73"),
   113 => (x"c3",x"87",x"ce",x"05"),
   114 => (x"de",x"ff",x"49",x"f4"),
   115 => (x"49",x"70",x"87",x"e8"),
   116 => (x"c2",x"02",x"99",x"c2"),
   117 => (x"73",x"4c",x"fa",x"87"),
   118 => (x"05",x"99",x"c8",x"49"),
   119 => (x"f5",x"c3",x"87",x"ce"),
   120 => (x"d1",x"de",x"ff",x"49"),
   121 => (x"c2",x"49",x"70",x"87"),
   122 => (x"87",x"d5",x"02",x"99"),
   123 => (x"bf",x"f9",x"e6",x"c2"),
   124 => (x"48",x"87",x"ca",x"02"),
   125 => (x"e6",x"c2",x"88",x"c1"),
   126 => (x"c2",x"c0",x"58",x"fd"),
   127 => (x"c1",x"4c",x"ff",x"87"),
   128 => (x"c4",x"49",x"73",x"4d"),
   129 => (x"87",x"ce",x"05",x"99"),
   130 => (x"ff",x"49",x"f2",x"c3"),
   131 => (x"70",x"87",x"e7",x"dd"),
   132 => (x"02",x"99",x"c2",x"49"),
   133 => (x"e6",x"c2",x"87",x"dc"),
   134 => (x"48",x"7e",x"bf",x"f9"),
   135 => (x"03",x"a8",x"b7",x"c7"),
   136 => (x"6e",x"87",x"cb",x"c0"),
   137 => (x"c2",x"80",x"c1",x"48"),
   138 => (x"c0",x"58",x"fd",x"e6"),
   139 => (x"4c",x"fe",x"87",x"c2"),
   140 => (x"fd",x"c3",x"4d",x"c1"),
   141 => (x"fd",x"dc",x"ff",x"49"),
   142 => (x"c2",x"49",x"70",x"87"),
   143 => (x"d5",x"c0",x"02",x"99"),
   144 => (x"f9",x"e6",x"c2",x"87"),
   145 => (x"c9",x"c0",x"02",x"bf"),
   146 => (x"f9",x"e6",x"c2",x"87"),
   147 => (x"c0",x"78",x"c0",x"48"),
   148 => (x"4c",x"fd",x"87",x"c2"),
   149 => (x"fa",x"c3",x"4d",x"c1"),
   150 => (x"d9",x"dc",x"ff",x"49"),
   151 => (x"c2",x"49",x"70",x"87"),
   152 => (x"d9",x"c0",x"02",x"99"),
   153 => (x"f9",x"e6",x"c2",x"87"),
   154 => (x"b7",x"c7",x"48",x"bf"),
   155 => (x"c9",x"c0",x"03",x"a8"),
   156 => (x"f9",x"e6",x"c2",x"87"),
   157 => (x"c0",x"78",x"c7",x"48"),
   158 => (x"4c",x"fc",x"87",x"c2"),
   159 => (x"b7",x"c0",x"4d",x"c1"),
   160 => (x"d1",x"c0",x"03",x"ac"),
   161 => (x"4a",x"66",x"c4",x"87"),
   162 => (x"6a",x"82",x"d8",x"c1"),
   163 => (x"87",x"c6",x"c0",x"02"),
   164 => (x"49",x"74",x"4b",x"6a"),
   165 => (x"1e",x"c0",x"0f",x"73"),
   166 => (x"c1",x"1e",x"f0",x"c3"),
   167 => (x"e4",x"f6",x"49",x"da"),
   168 => (x"70",x"86",x"c8",x"87"),
   169 => (x"e2",x"c0",x"02",x"98"),
   170 => (x"48",x"a6",x"c8",x"87"),
   171 => (x"bf",x"f9",x"e6",x"c2"),
   172 => (x"49",x"66",x"c8",x"78"),
   173 => (x"66",x"c4",x"91",x"cb"),
   174 => (x"70",x"80",x"71",x"48"),
   175 => (x"02",x"bf",x"6e",x"7e"),
   176 => (x"6e",x"87",x"c8",x"c0"),
   177 => (x"66",x"c8",x"4b",x"bf"),
   178 => (x"75",x"0f",x"73",x"49"),
   179 => (x"c8",x"c0",x"02",x"9d"),
   180 => (x"f9",x"e6",x"c2",x"87"),
   181 => (x"cd",x"f1",x"49",x"bf"),
   182 => (x"dc",x"cd",x"c2",x"87"),
   183 => (x"dd",x"c0",x"02",x"bf"),
   184 => (x"c7",x"c2",x"49",x"87"),
   185 => (x"02",x"98",x"70",x"87"),
   186 => (x"c2",x"87",x"d3",x"c0"),
   187 => (x"49",x"bf",x"f9",x"e6"),
   188 => (x"c0",x"87",x"f3",x"f0"),
   189 => (x"87",x"d3",x"f2",x"49"),
   190 => (x"48",x"dc",x"cd",x"c2"),
   191 => (x"8e",x"f4",x"78",x"c0"),
   192 => (x"0e",x"87",x"ed",x"f1"),
   193 => (x"5d",x"5c",x"5b",x"5e"),
   194 => (x"4c",x"71",x"1e",x"0e"),
   195 => (x"bf",x"f5",x"e6",x"c2"),
   196 => (x"a1",x"cd",x"c1",x"49"),
   197 => (x"81",x"d1",x"c1",x"4d"),
   198 => (x"9c",x"74",x"7e",x"69"),
   199 => (x"c4",x"87",x"cf",x"02"),
   200 => (x"7b",x"74",x"4b",x"a5"),
   201 => (x"bf",x"f5",x"e6",x"c2"),
   202 => (x"87",x"cc",x"f1",x"49"),
   203 => (x"9c",x"74",x"7b",x"6e"),
   204 => (x"c0",x"87",x"c4",x"05"),
   205 => (x"c1",x"87",x"c2",x"4b"),
   206 => (x"f1",x"49",x"73",x"4b"),
   207 => (x"66",x"d4",x"87",x"cd"),
   208 => (x"49",x"87",x"c7",x"02"),
   209 => (x"4a",x"70",x"87",x"da"),
   210 => (x"4a",x"c0",x"87",x"c2"),
   211 => (x"5a",x"e0",x"cd",x"c2"),
   212 => (x"87",x"dc",x"f0",x"26"),
   213 => (x"00",x"00",x"00",x"00"),
   214 => (x"00",x"00",x"00",x"00"),
   215 => (x"00",x"00",x"00",x"00"),
   216 => (x"ff",x"4a",x"71",x"1e"),
   217 => (x"72",x"49",x"bf",x"c8"),
   218 => (x"4f",x"26",x"48",x"a1"),
   219 => (x"bf",x"c8",x"ff",x"1e"),
   220 => (x"c0",x"c0",x"fe",x"89"),
   221 => (x"a9",x"c0",x"c0",x"c0"),
   222 => (x"c0",x"87",x"c4",x"01"),
   223 => (x"c1",x"87",x"c2",x"4a"),
   224 => (x"26",x"48",x"72",x"4a"),
   225 => (x"ce",x"c2",x"1e",x"4f"),
   226 => (x"c1",x"49",x"bf",x"ee"),
   227 => (x"f2",x"ce",x"c2",x"b9"),
   228 => (x"48",x"d4",x"ff",x"59"),
   229 => (x"ff",x"78",x"ff",x"c3"),
   230 => (x"e1",x"c0",x"48",x"d0"),
   231 => (x"48",x"d4",x"ff",x"78"),
   232 => (x"31",x"c4",x"78",x"c1"),
   233 => (x"d0",x"ff",x"78",x"71"),
   234 => (x"78",x"e0",x"c0",x"48"),
   235 => (x"00",x"00",x"4f",x"26"),
   236 => (x"5e",x"0e",x"00",x"00"),
   237 => (x"0e",x"5d",x"5c",x"5b"),
   238 => (x"bf",x"ec",x"4d",x"71"),
   239 => (x"ff",x"49",x"c5",x"4b"),
   240 => (x"70",x"87",x"f3",x"d6"),
   241 => (x"87",x"c7",x"05",x"98"),
   242 => (x"99",x"c2",x"49",x"73"),
   243 => (x"c2",x"87",x"c7",x"02"),
   244 => (x"c2",x"48",x"ed",x"d4"),
   245 => (x"49",x"c6",x"78",x"c0"),
   246 => (x"87",x"da",x"d6",x"ff"),
   247 => (x"c7",x"05",x"98",x"70"),
   248 => (x"c4",x"49",x"73",x"87"),
   249 => (x"87",x"c7",x"02",x"99"),
   250 => (x"48",x"ed",x"d4",x"c2"),
   251 => (x"c4",x"78",x"f0",x"c0"),
   252 => (x"c1",x"d6",x"ff",x"49"),
   253 => (x"05",x"98",x"70",x"87"),
   254 => (x"49",x"73",x"87",x"c7"),
   255 => (x"c6",x"02",x"99",x"c8"),
   256 => (x"ed",x"d4",x"c2",x"87"),
   257 => (x"cc",x"78",x"cc",x"48"),
   258 => (x"e9",x"d5",x"ff",x"49"),
   259 => (x"05",x"98",x"70",x"87"),
   260 => (x"49",x"73",x"87",x"c7"),
   261 => (x"c6",x"02",x"99",x"d0"),
   262 => (x"ed",x"d4",x"c2",x"87"),
   263 => (x"d0",x"78",x"c8",x"48"),
   264 => (x"49",x"75",x"1e",x"66"),
   265 => (x"87",x"f1",x"d7",x"ff"),
   266 => (x"bf",x"ed",x"d4",x"c2"),
   267 => (x"1e",x"66",x"d8",x"1e"),
   268 => (x"93",x"c2",x"4b",x"75"),
   269 => (x"94",x"c8",x"4c",x"75"),
   270 => (x"84",x"fd",x"e6",x"c2"),
   271 => (x"c4",x"ee",x"49",x"6c"),
   272 => (x"c2",x"7c",x"70",x"87"),
   273 => (x"1e",x"bf",x"ed",x"d4"),
   274 => (x"49",x"66",x"e0",x"c0"),
   275 => (x"71",x"29",x"b7",x"c2"),
   276 => (x"c2",x"93",x"c4",x"1e"),
   277 => (x"6b",x"83",x"c1",x"e7"),
   278 => (x"87",x"e9",x"ed",x"49"),
   279 => (x"e6",x"c2",x"7b",x"70"),
   280 => (x"49",x"75",x"1e",x"fd"),
   281 => (x"87",x"ce",x"d7",x"ff"),
   282 => (x"4d",x"26",x"8e",x"e8"),
   283 => (x"4b",x"26",x"4c",x"26"),
   284 => (x"73",x"1e",x"4f",x"26"),
   285 => (x"df",x"dc",x"c1",x"1e"),
   286 => (x"c2",x"50",x"c0",x"48"),
   287 => (x"c2",x"48",x"f0",x"d4"),
   288 => (x"c2",x"78",x"c0",x"c0"),
   289 => (x"48",x"bf",x"d4",x"e6"),
   290 => (x"e6",x"c2",x"b0",x"c1"),
   291 => (x"d7",x"ff",x"58",x"d8"),
   292 => (x"d3",x"c2",x"87",x"d4"),
   293 => (x"e3",x"fe",x"49",x"ee"),
   294 => (x"4b",x"70",x"87",x"c2"),
   295 => (x"bf",x"d4",x"e6",x"c2"),
   296 => (x"c2",x"98",x"fe",x"48"),
   297 => (x"ff",x"58",x"d8",x"e6"),
   298 => (x"73",x"87",x"fb",x"d6"),
   299 => (x"87",x"c7",x"05",x"9b"),
   300 => (x"48",x"fa",x"d3",x"c2"),
   301 => (x"c2",x"87",x"f4",x"c0"),
   302 => (x"48",x"bf",x"d4",x"e6"),
   303 => (x"e6",x"c2",x"b0",x"c1"),
   304 => (x"d6",x"ff",x"58",x"d8"),
   305 => (x"d4",x"c2",x"87",x"e0"),
   306 => (x"78",x"c1",x"48",x"f0"),
   307 => (x"48",x"df",x"dc",x"c1"),
   308 => (x"d4",x"c2",x"50",x"c1"),
   309 => (x"e2",x"fe",x"49",x"d1"),
   310 => (x"e6",x"c2",x"87",x"c2"),
   311 => (x"fe",x"48",x"bf",x"d4"),
   312 => (x"d8",x"e6",x"c2",x"98"),
   313 => (x"fd",x"d5",x"ff",x"58"),
   314 => (x"fe",x"48",x"c0",x"87"),
   315 => (x"45",x"56",x"87",x"c0"),
   316 => (x"45",x"52",x"54",x"43"),
   317 => (x"49",x"42",x"20",x"58"),
   318 => (x"45",x"56",x"00",x"4e"),
   319 => (x"45",x"52",x"54",x"43"),
   320 => (x"49",x"42",x"2e",x"58"),
   321 => (x"6f",x"6e",x"20",x"4e"),
   322 => (x"6f",x"66",x"20",x"74"),
   323 => (x"21",x"64",x"6e",x"75"),
   324 => (x"54",x"55",x"41",x"00"),
   325 => (x"4f",x"4f",x"42",x"4f"),
   326 => (x"43",x"45",x"56",x"54"),
   327 => (x"14",x"12",x"58",x"00"),
   328 => (x"1c",x"1b",x"1d",x"11"),
   329 => (x"49",x"4a",x"59",x"23"),
   330 => (x"eb",x"f2",x"f5",x"41"),
   331 => (x"00",x"00",x"80",x"f4"),
   332 => (x"00",x"00",x"80",x"00"),
		others => (others => x"00")
	);
	signal q1_local : word_t;

	-- Altera Quartus attributes
	attribute ramstyle: string;
	attribute ramstyle of ram: signal is "no_rw_check";

begin  -- rtl

	addr1 <= to_integer(unsigned(addr(ADDR_WIDTH-1 downto 0)));

	-- Reorganize the read data from the RAM to match the output
	q(7 downto 0) <= q1_local(3);
	q(15 downto 8) <= q1_local(2);
	q(23 downto 16) <= q1_local(1);
	q(31 downto 24) <= q1_local(0);

	process(clk)
	begin
		if(rising_edge(clk)) then 
			if(we = '1') then
				-- edit this code if using other than four bytes per word
				if (bytesel(3) = '1') then
					ram(addr1)(3) <= d(7 downto 0);
				end if;
				if (bytesel(2) = '1') then
					ram(addr1)(2) <= d(15 downto 8);
				end if;
				if (bytesel(1) = '1') then
					ram(addr1)(1) <= d(23 downto 16);
				end if;
				if (bytesel(0) = '1') then
					ram(addr1)(0) <= d(31 downto 24);
				end if;
			end if;
			q1_local <= ram(addr1);
		end if;
	end process;
  
end rtl;

