library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity controller_rom is
generic	(
	ADDR_WIDTH : integer := 8; -- ROM's address width (words, not bytes)
	COL_WIDTH  : integer := 8;  -- Column width (8bit -> byte)
	NB_COL     : integer := 4  -- Number of columns in memory
	);
port (
	clk : in std_logic;
	reset_n : in std_logic := '1';
	addr : in std_logic_vector(ADDR_WIDTH-1 downto 0);
	q : out std_logic_vector(31 downto 0);
	-- Allow writes - defaults supplied to simplify projects that don't need to write.
	d : in std_logic_vector(31 downto 0) := X"00000000";
	we : in std_logic := '0';
	bytesel : in std_logic_vector(3 downto 0) := "1111"
);
end entity;

architecture arch of controller_rom is

-- type word_t is std_logic_vector(31 downto 0);
type ram_type is array (0 to 2 ** ADDR_WIDTH - 1) of std_logic_vector(NB_COL * COL_WIDTH - 1 downto 0);

signal ram : ram_type :=
(

     0 => x"0487da01",
     1 => x"580e87dd",
     2 => x"0e5a595e",
     3 => x"00002927",
     4 => x"4a260f00",
     5 => x"48264926",
     6 => x"082680ff",
     7 => x"002d274f",
     8 => x"274f0000",
     9 => x"0000002a",
    10 => x"fd004f4f",
    11 => x"d0e7c287",
    12 => x"86c0c54e",
    13 => x"49d0e7c2",
    14 => x"48f4d4c2",
    15 => x"4040c089",
    16 => x"89d04040",
    17 => x"c187f603",
    18 => x"0087feda",
    19 => x"1e87fc98",
    20 => x"1e731e72",
    21 => x"02114812",
    22 => x"c34b87ca",
    23 => x"739b98df",
    24 => x"87f00288",
    25 => x"4a264b26",
    26 => x"731e4f26",
    27 => x"c11e721e",
    28 => x"87ca048b",
    29 => x"02114812",
    30 => x"028887c4",
    31 => x"4a2687f1",
    32 => x"4f264b26",
    33 => x"731e741e",
    34 => x"c11e721e",
    35 => x"87d0048b",
    36 => x"02114812",
    37 => x"c34c87ca",
    38 => x"749c98df",
    39 => x"87eb0288",
    40 => x"4b264a26",
    41 => x"4f264c26",
    42 => x"8148731e",
    43 => x"c502a973",
    44 => x"05531287",
    45 => x"4f2687f6",
    46 => x"4a66c41e",
    47 => x"51124871",
    48 => x"2687fb05",
    49 => x"4a711e4f",
    50 => x"484966c4",
    51 => x"a6c888c1",
    52 => x"02997158",
    53 => x"d4ff87d6",
    54 => x"78ffc348",
    55 => x"66c45268",
    56 => x"88c14849",
    57 => x"7158a6c8",
    58 => x"87ea0599",
    59 => x"731e4f26",
    60 => x"4bd4ff1e",
    61 => x"6b7bffc3",
    62 => x"7bffc34a",
    63 => x"32c8496b",
    64 => x"ffc3b172",
    65 => x"c84a6b7b",
    66 => x"c3b27131",
    67 => x"496b7bff",
    68 => x"b17232c8",
    69 => x"87c44871",
    70 => x"4c264d26",
    71 => x"4f264b26",
    72 => x"5c5b5e0e",
    73 => x"4a710e5d",
    74 => x"724cd4ff",
    75 => x"99ffc349",
    76 => x"d4c27c71",
    77 => x"c805bff4",
    78 => x"4866d087",
    79 => x"a6d430c9",
    80 => x"4966d058",
    81 => x"ffc329d8",
    82 => x"d07c7199",
    83 => x"29d04966",
    84 => x"7199ffc3",
    85 => x"4966d07c",
    86 => x"ffc329c8",
    87 => x"d07c7199",
    88 => x"ffc34966",
    89 => x"727c7199",
    90 => x"c329d049",
    91 => x"7c7199ff",
    92 => x"f0c94b6c",
    93 => x"ffc34dff",
    94 => x"87d005ab",
    95 => x"6c7cffc3",
    96 => x"028dc14b",
    97 => x"ffc387c6",
    98 => x"87f002ab",
    99 => x"c7fe4873",
   100 => x"49c01e87",
   101 => x"c348d4ff",
   102 => x"81c178ff",
   103 => x"a9b7c8c3",
   104 => x"2687f104",
   105 => x"1e731e4f",
   106 => x"f8c487e7",
   107 => x"1ec04bdf",
   108 => x"c1f0ffc0",
   109 => x"e7fd49f7",
   110 => x"c186c487",
   111 => x"eac005a8",
   112 => x"48d4ff87",
   113 => x"c178ffc3",
   114 => x"c0c0c0c0",
   115 => x"e1c01ec0",
   116 => x"49e9c1f0",
   117 => x"c487c9fd",
   118 => x"05987086",
   119 => x"d4ff87ca",
   120 => x"78ffc348",
   121 => x"87cb48c1",
   122 => x"c187e6fe",
   123 => x"fdfe058b",
   124 => x"fc48c087",
   125 => x"731e87e6",
   126 => x"48d4ff1e",
   127 => x"d378ffc3",
   128 => x"c01ec04b",
   129 => x"c1c1f0ff",
   130 => x"87d4fc49",
   131 => x"987086c4",
   132 => x"ff87ca05",
   133 => x"ffc348d4",
   134 => x"cb48c178",
   135 => x"87f1fd87",
   136 => x"ff058bc1",
   137 => x"48c087db",
   138 => x"0e87f1fb",
   139 => x"0e5c5b5e",
   140 => x"fd4cd4ff",
   141 => x"eac687db",
   142 => x"f0e1c01e",
   143 => x"fb49c8c1",
   144 => x"86c487de",
   145 => x"c802a8c1",
   146 => x"87eafe87",
   147 => x"e2c148c0",
   148 => x"87dafa87",
   149 => x"ffcf4970",
   150 => x"eac699ff",
   151 => x"87c802a9",
   152 => x"c087d3fe",
   153 => x"87cbc148",
   154 => x"c07cffc3",
   155 => x"f4fc4bf1",
   156 => x"02987087",
   157 => x"c087ebc0",
   158 => x"f0ffc01e",
   159 => x"fa49fac1",
   160 => x"86c487de",
   161 => x"d9059870",
   162 => x"7cffc387",
   163 => x"ffc3496c",
   164 => x"7c7c7c7c",
   165 => x"0299c0c1",
   166 => x"48c187c4",
   167 => x"48c087d5",
   168 => x"abc287d1",
   169 => x"c087c405",
   170 => x"c187c848",
   171 => x"fdfe058b",
   172 => x"f948c087",
   173 => x"731e87e4",
   174 => x"f4d4c21e",
   175 => x"c778c148",
   176 => x"48d0ff4b",
   177 => x"c8fb78c2",
   178 => x"48d0ff87",
   179 => x"1ec078c3",
   180 => x"c1d0e5c0",
   181 => x"c7f949c0",
   182 => x"c186c487",
   183 => x"87c105a8",
   184 => x"05abc24b",
   185 => x"48c087c5",
   186 => x"c187f9c0",
   187 => x"d0ff058b",
   188 => x"87f7fc87",
   189 => x"58f8d4c2",
   190 => x"cd059870",
   191 => x"c01ec187",
   192 => x"d0c1f0ff",
   193 => x"87d8f849",
   194 => x"d4ff86c4",
   195 => x"78ffc348",
   196 => x"c287fcc2",
   197 => x"ff58fcd4",
   198 => x"78c248d0",
   199 => x"c348d4ff",
   200 => x"48c178ff",
   201 => x"0e87f5f7",
   202 => x"5d5c5b5e",
   203 => x"c04b710e",
   204 => x"cdeec54c",
   205 => x"d4ff4adf",
   206 => x"78ffc348",
   207 => x"fec34968",
   208 => x"fdc005a9",
   209 => x"734d7087",
   210 => x"87cc029b",
   211 => x"731e66d0",
   212 => x"87f1f549",
   213 => x"87d686c4",
   214 => x"c448d0ff",
   215 => x"ffc378d1",
   216 => x"4866d07d",
   217 => x"a6d488c1",
   218 => x"05987058",
   219 => x"d4ff87f0",
   220 => x"78ffc348",
   221 => x"059b7378",
   222 => x"d0ff87c5",
   223 => x"c178d048",
   224 => x"8ac14c4a",
   225 => x"87eefe05",
   226 => x"cbf64874",
   227 => x"1e731e87",
   228 => x"4bc04a71",
   229 => x"c348d4ff",
   230 => x"d0ff78ff",
   231 => x"78c3c448",
   232 => x"c348d4ff",
   233 => x"1e7278ff",
   234 => x"c1f0ffc0",
   235 => x"eff549d1",
   236 => x"7086c487",
   237 => x"87d20598",
   238 => x"cc1ec0c8",
   239 => x"e6fd4966",
   240 => x"7086c487",
   241 => x"48d0ff4b",
   242 => x"487378c2",
   243 => x"0e87cdf5",
   244 => x"5d5c5b5e",
   245 => x"c01ec00e",
   246 => x"c9c1f0ff",
   247 => x"87c0f549",
   248 => x"d4c21ed2",
   249 => x"fefc49fc",
   250 => x"c086c887",
   251 => x"d284c14c",
   252 => x"f804acb7",
   253 => x"fcd4c287",
   254 => x"c349bf97",
   255 => x"c0c199c0",
   256 => x"e7c005a9",
   257 => x"c3d5c287",
   258 => x"d049bf97",
   259 => x"c4d5c231",
   260 => x"c84abf97",
   261 => x"c2b17232",
   262 => x"bf97c5d5",
   263 => x"4c71b14a",
   264 => x"ffffffcf",
   265 => x"ca84c19c",
   266 => x"87e7c134",
   267 => x"97c5d5c2",
   268 => x"31c149bf",
   269 => x"d5c299c6",
   270 => x"4abf97c6",
   271 => x"722ab7c7",
   272 => x"c1d5c2b1",
   273 => x"4d4abf97",
   274 => x"d5c29dcf",
   275 => x"4abf97c2",
   276 => x"32ca9ac3",
   277 => x"97c3d5c2",
   278 => x"33c24bbf",
   279 => x"d5c2b273",
   280 => x"4bbf97c4",
   281 => x"c69bc0c3",
   282 => x"b2732bb7",
   283 => x"48c181c2",
   284 => x"49703071",
   285 => x"307548c1",
   286 => x"4c724d70",
   287 => x"947184c1",
   288 => x"adb7c0c8",
   289 => x"c187cc06",
   290 => x"c82db734",
   291 => x"01adb7c0",
   292 => x"7487f4ff",
   293 => x"87c0f248",
   294 => x"5c5b5e0e",
   295 => x"86f80e5d",
   296 => x"48e2ddc2",
   297 => x"d5c278c0",
   298 => x"49c01eda",
   299 => x"c487defb",
   300 => x"05987086",
   301 => x"48c087c5",
   302 => x"c087cec9",
   303 => x"c07ec14d",
   304 => x"49bfc1ee",
   305 => x"4ad0d6c2",
   306 => x"ee4bc871",
   307 => x"987087dc",
   308 => x"c087c205",
   309 => x"fdedc07e",
   310 => x"d6c249bf",
   311 => x"c8714aec",
   312 => x"87c6ee4b",
   313 => x"c2059870",
   314 => x"6e7ec087",
   315 => x"87fdc002",
   316 => x"bfe0dcc2",
   317 => x"d8ddc24d",
   318 => x"487ebf9f",
   319 => x"a8ead6c5",
   320 => x"c287c705",
   321 => x"4dbfe0dc",
   322 => x"486e87ce",
   323 => x"a8d5e9ca",
   324 => x"c087c502",
   325 => x"87f1c748",
   326 => x"1edad5c2",
   327 => x"ecf94975",
   328 => x"7086c487",
   329 => x"87c50598",
   330 => x"dcc748c0",
   331 => x"fdedc087",
   332 => x"d6c249bf",
   333 => x"c8714aec",
   334 => x"87eeec4b",
   335 => x"c8059870",
   336 => x"e2ddc287",
   337 => x"da78c148",
   338 => x"c1eec087",
   339 => x"d6c249bf",
   340 => x"c8714ad0",
   341 => x"87d2ec4b",
   342 => x"c0029870",
   343 => x"48c087c5",
   344 => x"c287e6c6",
   345 => x"bf97d8dd",
   346 => x"a9d5c149",
   347 => x"87cdc005",
   348 => x"97d9ddc2",
   349 => x"eac249bf",
   350 => x"c5c002a9",
   351 => x"c648c087",
   352 => x"d5c287c7",
   353 => x"7ebf97da",
   354 => x"a8e9c348",
   355 => x"87cec002",
   356 => x"ebc3486e",
   357 => x"c5c002a8",
   358 => x"c548c087",
   359 => x"d5c287eb",
   360 => x"49bf97e5",
   361 => x"ccc00599",
   362 => x"e6d5c287",
   363 => x"c249bf97",
   364 => x"c5c002a9",
   365 => x"c548c087",
   366 => x"d5c287cf",
   367 => x"48bf97e7",
   368 => x"58deddc2",
   369 => x"c1484c70",
   370 => x"e2ddc288",
   371 => x"e8d5c258",
   372 => x"7549bf97",
   373 => x"e9d5c281",
   374 => x"c84abf97",
   375 => x"7ea17232",
   376 => x"48efe1c2",
   377 => x"d5c2786e",
   378 => x"48bf97ea",
   379 => x"c258a6c8",
   380 => x"02bfe2dd",
   381 => x"c087d4c2",
   382 => x"49bffded",
   383 => x"4aecd6c2",
   384 => x"e94bc871",
   385 => x"987087e4",
   386 => x"87c5c002",
   387 => x"f8c348c0",
   388 => x"daddc287",
   389 => x"e2c24cbf",
   390 => x"d5c25cc3",
   391 => x"49bf97ff",
   392 => x"d5c231c8",
   393 => x"4abf97fe",
   394 => x"d6c249a1",
   395 => x"4abf97c0",
   396 => x"a17232d0",
   397 => x"c1d6c249",
   398 => x"d84abf97",
   399 => x"49a17232",
   400 => x"c29166c4",
   401 => x"81bfefe1",
   402 => x"59f7e1c2",
   403 => x"97c7d6c2",
   404 => x"32c84abf",
   405 => x"97c6d6c2",
   406 => x"4aa24bbf",
   407 => x"97c8d6c2",
   408 => x"33d04bbf",
   409 => x"c24aa273",
   410 => x"bf97c9d6",
   411 => x"d89bcf4b",
   412 => x"4aa27333",
   413 => x"5afbe1c2",
   414 => x"bff7e1c2",
   415 => x"748ac24a",
   416 => x"fbe1c292",
   417 => x"78a17248",
   418 => x"c287cac1",
   419 => x"bf97ecd5",
   420 => x"c231c849",
   421 => x"bf97ebd5",
   422 => x"c249a14a",
   423 => x"c259eadd",
   424 => x"49bfe6dd",
   425 => x"ffc731c5",
   426 => x"c229c981",
   427 => x"c259c3e2",
   428 => x"bf97f1d5",
   429 => x"c232c84a",
   430 => x"bf97f0d5",
   431 => x"c44aa24b",
   432 => x"826e9266",
   433 => x"5affe1c2",
   434 => x"48f7e1c2",
   435 => x"e1c278c0",
   436 => x"a17248f3",
   437 => x"c3e2c278",
   438 => x"f7e1c248",
   439 => x"e2c278bf",
   440 => x"e1c248c7",
   441 => x"c278bffb",
   442 => x"02bfe2dd",
   443 => x"7487c9c0",
   444 => x"7030c448",
   445 => x"87c9c07e",
   446 => x"bfffe1c2",
   447 => x"7030c448",
   448 => x"e6ddc27e",
   449 => x"c1786e48",
   450 => x"268ef848",
   451 => x"264c264d",
   452 => x"0e4f264b",
   453 => x"5d5c5b5e",
   454 => x"c24a710e",
   455 => x"02bfe2dd",
   456 => x"4b7287cb",
   457 => x"4c722bc7",
   458 => x"c99cffc1",
   459 => x"c84b7287",
   460 => x"c34c722b",
   461 => x"e1c29cff",
   462 => x"c083bfef",
   463 => x"abbff9ed",
   464 => x"c087d902",
   465 => x"c25bfded",
   466 => x"731edad5",
   467 => x"87fdf049",
   468 => x"987086c4",
   469 => x"c087c505",
   470 => x"87e6c048",
   471 => x"bfe2ddc2",
   472 => x"7487d202",
   473 => x"c291c449",
   474 => x"6981dad5",
   475 => x"ffffcf4d",
   476 => x"cb9dffff",
   477 => x"c2497487",
   478 => x"dad5c291",
   479 => x"4d699f81",
   480 => x"c6fe4875",
   481 => x"5b5e0e87",
   482 => x"1e0e5d5c",
   483 => x"1ec04d71",
   484 => x"c9c849c1",
   485 => x"7086c487",
   486 => x"c1029c4c",
   487 => x"ddc287c0",
   488 => x"49754aea",
   489 => x"7087e8e2",
   490 => x"f1c00298",
   491 => x"754a7487",
   492 => x"e34bcb49",
   493 => x"987087ce",
   494 => x"87e2c002",
   495 => x"9c741ec0",
   496 => x"c487c702",
   497 => x"78c048a6",
   498 => x"a6c487c5",
   499 => x"c478c148",
   500 => x"c9c74966",
   501 => x"7086c487",
   502 => x"ff059c4c",
   503 => x"487487c0",
   504 => x"87e7fc26",
   505 => x"5c5b5e0e",
   506 => x"711e0e5d",
   507 => x"c5059b4b",
   508 => x"c148c087",
   509 => x"a3c887e5",
   510 => x"d47dc04d",
   511 => x"87c70266",
   512 => x"bf9766d4",
   513 => x"c087c505",
   514 => x"87cfc148",
   515 => x"fd4966d4",
   516 => x"4c7087f3",
   517 => x"c0c1029c",
   518 => x"49a4dc87",
   519 => x"a4da7d69",
   520 => x"4aa3c449",
   521 => x"c27a699f",
   522 => x"02bfe2dd",
   523 => x"a4d487d2",
   524 => x"49699f49",
   525 => x"99ffffc0",
   526 => x"30d04871",
   527 => x"87c27e70",
   528 => x"496e7ec0",
   529 => x"70806a48",
   530 => x"cc7bc07a",
   531 => x"796a49a3",
   532 => x"c049a3d0",
   533 => x"c248c179",
   534 => x"2648c087",
   535 => x"0e87ecfa",
   536 => x"5d5c5b5e",
   537 => x"9c4c710e",
   538 => x"87cac102",
   539 => x"6949a4c8",
   540 => x"87c2c102",
   541 => x"6c4a66d0",
   542 => x"a6d48249",
   543 => x"4d66d05a",
   544 => x"deddc2b9",
   545 => x"baff4abf",
   546 => x"99719972",
   547 => x"87e4c002",
   548 => x"6b4ba4c4",
   549 => x"87fbf949",
   550 => x"ddc27b70",
   551 => x"6c49bfda",
   552 => x"757c7181",
   553 => x"deddc2b9",
   554 => x"baff4abf",
   555 => x"99719972",
   556 => x"87dcff05",
   557 => x"d2f97c75",
   558 => x"1e731e87",
   559 => x"029b4b71",
   560 => x"a3c887c7",
   561 => x"c5056949",
   562 => x"c048c087",
   563 => x"e1c287f7",
   564 => x"c44abff3",
   565 => x"496949a3",
   566 => x"ddc289c2",
   567 => x"7191bfda",
   568 => x"ddc24aa2",
   569 => x"6b49bfde",
   570 => x"4aa27199",
   571 => x"5afdedc0",
   572 => x"721e66c8",
   573 => x"87d5ea49",
   574 => x"987086c4",
   575 => x"c087c405",
   576 => x"c187c248",
   577 => x"87c7f848",
   578 => x"711e731e",
   579 => x"c0029b4b",
   580 => x"e2c287e4",
   581 => x"4a735bc7",
   582 => x"ddc28ac2",
   583 => x"9249bfda",
   584 => x"bff3e1c2",
   585 => x"c2807248",
   586 => x"7158cbe2",
   587 => x"c230c448",
   588 => x"c058eadd",
   589 => x"e2c287ed",
   590 => x"e1c248c3",
   591 => x"c278bff7",
   592 => x"c248c7e2",
   593 => x"78bffbe1",
   594 => x"bfe2ddc2",
   595 => x"c287c902",
   596 => x"49bfdadd",
   597 => x"87c731c4",
   598 => x"bfffe1c2",
   599 => x"c231c449",
   600 => x"f659eadd",
   601 => x"5e0e87e9",
   602 => x"710e5c5b",
   603 => x"724bc04a",
   604 => x"e1c0029a",
   605 => x"49a2da87",
   606 => x"c24b699f",
   607 => x"02bfe2dd",
   608 => x"a2d487cf",
   609 => x"49699f49",
   610 => x"ffffc04c",
   611 => x"c234d09c",
   612 => x"744cc087",
   613 => x"4973b349",
   614 => x"f587edfd",
   615 => x"5e0e87ef",
   616 => x"0e5d5c5b",
   617 => x"4a7186f4",
   618 => x"9a727ec0",
   619 => x"c287d802",
   620 => x"c048d6d5",
   621 => x"ced5c278",
   622 => x"c7e2c248",
   623 => x"d5c278bf",
   624 => x"e2c248d2",
   625 => x"c278bfc3",
   626 => x"c048f7dd",
   627 => x"e6ddc250",
   628 => x"d5c249bf",
   629 => x"714abfd6",
   630 => x"c9c403aa",
   631 => x"cf497287",
   632 => x"e9c00599",
   633 => x"f9edc087",
   634 => x"ced5c248",
   635 => x"d5c278bf",
   636 => x"d5c21eda",
   637 => x"c249bfce",
   638 => x"c148ced5",
   639 => x"e67178a1",
   640 => x"86c487cb",
   641 => x"48f5edc0",
   642 => x"78dad5c2",
   643 => x"edc087cc",
   644 => x"c048bff5",
   645 => x"edc080e0",
   646 => x"d5c258f9",
   647 => x"c148bfd6",
   648 => x"dad5c280",
   649 => x"0b752758",
   650 => x"97bf0000",
   651 => x"029d4dbf",
   652 => x"c387e3c2",
   653 => x"c202ade5",
   654 => x"edc087dc",
   655 => x"cb4bbff5",
   656 => x"4c1149a3",
   657 => x"c105accf",
   658 => x"497587d2",
   659 => x"89c199df",
   660 => x"ddc291cd",
   661 => x"a3c181ea",
   662 => x"c351124a",
   663 => x"51124aa3",
   664 => x"124aa3c5",
   665 => x"4aa3c751",
   666 => x"a3c95112",
   667 => x"ce51124a",
   668 => x"51124aa3",
   669 => x"124aa3d0",
   670 => x"4aa3d251",
   671 => x"a3d45112",
   672 => x"d651124a",
   673 => x"51124aa3",
   674 => x"124aa3d8",
   675 => x"4aa3dc51",
   676 => x"a3de5112",
   677 => x"c151124a",
   678 => x"87fac07e",
   679 => x"99c84974",
   680 => x"87ebc005",
   681 => x"99d04974",
   682 => x"dc87d105",
   683 => x"cbc00266",
   684 => x"dc497387",
   685 => x"98700f66",
   686 => x"87d3c002",
   687 => x"c6c0056e",
   688 => x"eaddc287",
   689 => x"c050c048",
   690 => x"48bff5ed",
   691 => x"c287e1c2",
   692 => x"c048f7dd",
   693 => x"ddc27e50",
   694 => x"c249bfe6",
   695 => x"4abfd6d5",
   696 => x"fb04aa71",
   697 => x"e2c287f7",
   698 => x"c005bfc7",
   699 => x"ddc287c8",
   700 => x"c102bfe2",
   701 => x"d5c287f8",
   702 => x"f049bfd2",
   703 => x"497087d5",
   704 => x"59d6d5c2",
   705 => x"c248a6c4",
   706 => x"78bfd2d5",
   707 => x"bfe2ddc2",
   708 => x"87d8c002",
   709 => x"cf4966c4",
   710 => x"f8ffffff",
   711 => x"c002a999",
   712 => x"4cc087c5",
   713 => x"c187e1c0",
   714 => x"87dcc04c",
   715 => x"cf4966c4",
   716 => x"a999f8ff",
   717 => x"87c8c002",
   718 => x"c048a6c8",
   719 => x"87c5c078",
   720 => x"c148a6c8",
   721 => x"4c66c878",
   722 => x"c0059c74",
   723 => x"66c487e0",
   724 => x"c289c249",
   725 => x"4abfdadd",
   726 => x"f3e1c291",
   727 => x"d5c24abf",
   728 => x"a17248ce",
   729 => x"d6d5c278",
   730 => x"f978c048",
   731 => x"48c087df",
   732 => x"d6ee8ef4",
   733 => x"00000087",
   734 => x"ffffff00",
   735 => x"000b85ff",
   736 => x"000b8e00",
   737 => x"54414600",
   738 => x"20203233",
   739 => x"41460020",
   740 => x"20363154",
   741 => x"1e002020",
   742 => x"c348d4ff",
   743 => x"486878ff",
   744 => x"ff1e4f26",
   745 => x"ffc348d4",
   746 => x"48d0ff78",
   747 => x"ff78e1c0",
   748 => x"78d448d4",
   749 => x"48cbe2c2",
   750 => x"50bfd4ff",
   751 => x"ff1e4f26",
   752 => x"e0c048d0",
   753 => x"1e4f2678",
   754 => x"7087ccff",
   755 => x"c6029949",
   756 => x"a9fbc087",
   757 => x"7187f105",
   758 => x"0e4f2648",
   759 => x"0e5c5b5e",
   760 => x"4cc04b71",
   761 => x"7087f0fe",
   762 => x"c0029949",
   763 => x"ecc087f9",
   764 => x"f2c002a9",
   765 => x"a9fbc087",
   766 => x"87ebc002",
   767 => x"acb766cc",
   768 => x"d087c703",
   769 => x"87c20266",
   770 => x"99715371",
   771 => x"c187c202",
   772 => x"87c3fe84",
   773 => x"02994970",
   774 => x"ecc087cd",
   775 => x"87c702a9",
   776 => x"05a9fbc0",
   777 => x"d087d5ff",
   778 => x"87c30266",
   779 => x"c07b97c0",
   780 => x"c405a9ec",
   781 => x"c54a7487",
   782 => x"c04a7487",
   783 => x"48728a0a",
   784 => x"4d2687c2",
   785 => x"4b264c26",
   786 => x"fd1e4f26",
   787 => x"497087c9",
   788 => x"a9b7f0c0",
   789 => x"c087ca04",
   790 => x"01a9b7f9",
   791 => x"f0c087c3",
   792 => x"b7c1c189",
   793 => x"87ca04a9",
   794 => x"a9b7dac1",
   795 => x"c087c301",
   796 => x"487189f7",
   797 => x"5e0e4f26",
   798 => x"710e5c5b",
   799 => x"4cd4ff4a",
   800 => x"e9c04972",
   801 => x"9b4b7087",
   802 => x"c187c202",
   803 => x"48d0ff8b",
   804 => x"d5c178c5",
   805 => x"c649737c",
   806 => x"dfdcc131",
   807 => x"484abf97",
   808 => x"7c70b071",
   809 => x"c448d0ff",
   810 => x"fe487378",
   811 => x"5e0e87d6",
   812 => x"0e5d5c5b",
   813 => x"4c7186f8",
   814 => x"e5fb7ec0",
   815 => x"c04bc087",
   816 => x"bf97dbf5",
   817 => x"04a9c049",
   818 => x"fafb87cf",
   819 => x"c083c187",
   820 => x"bf97dbf5",
   821 => x"f106ab49",
   822 => x"dbf5c087",
   823 => x"cf02bf97",
   824 => x"87f3fa87",
   825 => x"02994970",
   826 => x"ecc087c6",
   827 => x"87f105a9",
   828 => x"e2fa4bc0",
   829 => x"fa4d7087",
   830 => x"a6c887dd",
   831 => x"87d7fa58",
   832 => x"83c14a70",
   833 => x"9749a4c8",
   834 => x"02ad4969",
   835 => x"ffc087c7",
   836 => x"e7c005ad",
   837 => x"49a4c987",
   838 => x"c4496997",
   839 => x"c702a966",
   840 => x"ffc04887",
   841 => x"87d405a8",
   842 => x"9749a4ca",
   843 => x"02aa4969",
   844 => x"ffc087c6",
   845 => x"87c405aa",
   846 => x"87d07ec1",
   847 => x"02adecc0",
   848 => x"fbc087c6",
   849 => x"87c405ad",
   850 => x"7ec14bc0",
   851 => x"e1fe026e",
   852 => x"87eaf987",
   853 => x"8ef84873",
   854 => x"0087e7fb",
   855 => x"5c5b5e0e",
   856 => x"711e0e5d",
   857 => x"4bd4ff4d",
   858 => x"e2c21e75",
   859 => x"f3e949d0",
   860 => x"7086c487",
   861 => x"d5c30298",
   862 => x"d8e2c287",
   863 => x"49754cbf",
   864 => x"ff87f3fb",
   865 => x"78c548d0",
   866 => x"c07bd6c1",
   867 => x"49a2754a",
   868 => x"82c17b11",
   869 => x"04aab7cb",
   870 => x"4acc87f3",
   871 => x"c17bffc3",
   872 => x"b7e0c082",
   873 => x"87f404aa",
   874 => x"c448d0ff",
   875 => x"7bffc378",
   876 => x"d3c178c5",
   877 => x"c47bc17b",
   878 => x"029c7478",
   879 => x"c287ffc1",
   880 => x"c87edad5",
   881 => x"c08c4dc0",
   882 => x"c603acb7",
   883 => x"a4c0c887",
   884 => x"c84cc04d",
   885 => x"dc05adc0",
   886 => x"cbe2c287",
   887 => x"d049bf97",
   888 => x"87d10299",
   889 => x"e2c21ec0",
   890 => x"cceb49d0",
   891 => x"7086c487",
   892 => x"eec04a49",
   893 => x"dad5c287",
   894 => x"d0e2c21e",
   895 => x"87f9ea49",
   896 => x"497086c4",
   897 => x"48d0ff4a",
   898 => x"c178c5c8",
   899 => x"976e7bd4",
   900 => x"486e7bbf",
   901 => x"7e7080c1",
   902 => x"ff058dc1",
   903 => x"d0ff87f0",
   904 => x"7278c448",
   905 => x"87c5059a",
   906 => x"e3c048c0",
   907 => x"c21ec187",
   908 => x"e849d0e2",
   909 => x"86c487e9",
   910 => x"fe059c74",
   911 => x"d0ff87c1",
   912 => x"c178c548",
   913 => x"7bc07bd3",
   914 => x"48c178c4",
   915 => x"48c087c2",
   916 => x"264d2626",
   917 => x"264b264c",
   918 => x"5b5e0e4f",
   919 => x"1e0e5d5c",
   920 => x"4cc04b71",
   921 => x"c004ab4d",
   922 => x"f2c087e8",
   923 => x"9d751eee",
   924 => x"c087c402",
   925 => x"c187c24a",
   926 => x"ec49724a",
   927 => x"86c487e0",
   928 => x"84c17e70",
   929 => x"87c2056e",
   930 => x"85c14c73",
   931 => x"ff06ac73",
   932 => x"486e87d8",
   933 => x"87f9fe26",
   934 => x"c44a711e",
   935 => x"87c50566",
   936 => x"f7fa4972",
   937 => x"0e4f2687",
   938 => x"5d5c5b5e",
   939 => x"4c711e0e",
   940 => x"c291de49",
   941 => x"714df8e2",
   942 => x"026d9785",
   943 => x"c287dcc1",
   944 => x"4abfe4e2",
   945 => x"49728274",
   946 => x"7087cefe",
   947 => x"c0026e7e",
   948 => x"e2c287f2",
   949 => x"4a6e4bec",
   950 => x"c7ff49cb",
   951 => x"4b7487ca",
   952 => x"dcc193cb",
   953 => x"83c483ef",
   954 => x"7bdffcc0",
   955 => x"c0c14974",
   956 => x"7b7587f4",
   957 => x"97e0dcc1",
   958 => x"c21e49bf",
   959 => x"fe49ece2",
   960 => x"86c487d6",
   961 => x"c0c14974",
   962 => x"49c087dc",
   963 => x"87fbc1c1",
   964 => x"48cce2c2",
   965 => x"49c178c0",
   966 => x"2687c0dd",
   967 => x"4c87f2fc",
   968 => x"6964616f",
   969 => x"2e2e676e",
   970 => x"5e0e002e",
   971 => x"710e5c5b",
   972 => x"e2c24a4b",
   973 => x"7282bfe4",
   974 => x"87ddfc49",
   975 => x"029c4c70",
   976 => x"e84987c4",
   977 => x"e2c287e0",
   978 => x"78c048e4",
   979 => x"cadc49c1",
   980 => x"87fffb87",
   981 => x"5c5b5e0e",
   982 => x"86f40e5d",
   983 => x"4ddad5c2",
   984 => x"a6c44cc0",
   985 => x"c278c048",
   986 => x"49bfe4e2",
   987 => x"c106a9c0",
   988 => x"d5c287c1",
   989 => x"029848da",
   990 => x"c087f8c0",
   991 => x"c81eeef2",
   992 => x"87c70266",
   993 => x"c048a6c4",
   994 => x"c487c578",
   995 => x"78c148a6",
   996 => x"e84966c4",
   997 => x"86c487c8",
   998 => x"84c14d70",
   999 => x"c14866c4",
  1000 => x"58a6c880",
  1001 => x"bfe4e2c2",
  1002 => x"c603ac49",
  1003 => x"059d7587",
  1004 => x"c087c8ff",
  1005 => x"029d754c",
  1006 => x"c087e0c3",
  1007 => x"c81eeef2",
  1008 => x"87c70266",
  1009 => x"c048a6cc",
  1010 => x"cc87c578",
  1011 => x"78c148a6",
  1012 => x"e74966cc",
  1013 => x"86c487c8",
  1014 => x"026e7e70",
  1015 => x"6e87e9c2",
  1016 => x"9781cb49",
  1017 => x"99d04969",
  1018 => x"87d6c102",
  1019 => x"4aeafcc0",
  1020 => x"91cb4974",
  1021 => x"81efdcc1",
  1022 => x"81c87972",
  1023 => x"7451ffc3",
  1024 => x"c291de49",
  1025 => x"714df8e2",
  1026 => x"97c1c285",
  1027 => x"49a5c17d",
  1028 => x"c251e0c0",
  1029 => x"bf97eadd",
  1030 => x"c187d202",
  1031 => x"4ba5c284",
  1032 => x"4aeaddc2",
  1033 => x"c1ff49db",
  1034 => x"dbc187fe",
  1035 => x"49a5cd87",
  1036 => x"84c151c0",
  1037 => x"6e4ba5c2",
  1038 => x"ff49cb4a",
  1039 => x"c187e9c1",
  1040 => x"fac087c6",
  1041 => x"49744ae7",
  1042 => x"dcc191cb",
  1043 => x"797281ef",
  1044 => x"97eaddc2",
  1045 => x"87d802bf",
  1046 => x"91de4974",
  1047 => x"e2c284c1",
  1048 => x"83714bf8",
  1049 => x"4aeaddc2",
  1050 => x"c0ff49dd",
  1051 => x"87d887fa",
  1052 => x"93de4b74",
  1053 => x"83f8e2c2",
  1054 => x"c049a3cb",
  1055 => x"7384c151",
  1056 => x"49cb4a6e",
  1057 => x"87e0c0ff",
  1058 => x"c14866c4",
  1059 => x"58a6c880",
  1060 => x"c003acc7",
  1061 => x"056e87c5",
  1062 => x"7487e0fc",
  1063 => x"f68ef448",
  1064 => x"731e87ef",
  1065 => x"494b711e",
  1066 => x"dcc191cb",
  1067 => x"a1c881ef",
  1068 => x"dfdcc14a",
  1069 => x"c9501248",
  1070 => x"f5c04aa1",
  1071 => x"501248db",
  1072 => x"dcc181ca",
  1073 => x"501148e0",
  1074 => x"97e0dcc1",
  1075 => x"c01e49bf",
  1076 => x"87c4f749",
  1077 => x"48cce2c2",
  1078 => x"49c178de",
  1079 => x"2687fcd5",
  1080 => x"1e87f2f5",
  1081 => x"cb494a71",
  1082 => x"efdcc191",
  1083 => x"1181c881",
  1084 => x"d0e2c248",
  1085 => x"e4e2c258",
  1086 => x"c178c048",
  1087 => x"87dbd549",
  1088 => x"c01e4f26",
  1089 => x"c2fac049",
  1090 => x"1e4f2687",
  1091 => x"d2029971",
  1092 => x"c4dec187",
  1093 => x"f750c048",
  1094 => x"e3c3c180",
  1095 => x"e8dcc140",
  1096 => x"c187ce78",
  1097 => x"c148c0de",
  1098 => x"fc78e1dc",
  1099 => x"c2c4c180",
  1100 => x"0e4f2678",
  1101 => x"0e5c5b5e",
  1102 => x"cb4a4c71",
  1103 => x"efdcc192",
  1104 => x"49a2c882",
  1105 => x"974ba2c9",
  1106 => x"971e4b6b",
  1107 => x"ca1e4969",
  1108 => x"c0491282",
  1109 => x"c087fde4",
  1110 => x"87ffd349",
  1111 => x"f7c04974",
  1112 => x"8ef887c4",
  1113 => x"1e87ecf3",
  1114 => x"4b711e73",
  1115 => x"87c3ff49",
  1116 => x"fefe4973",
  1117 => x"87ddf387",
  1118 => x"711e731e",
  1119 => x"4aa3c64b",
  1120 => x"c187db02",
  1121 => x"87d6028a",
  1122 => x"dac1028a",
  1123 => x"c0028a87",
  1124 => x"028a87fc",
  1125 => x"8a87e1c0",
  1126 => x"c187cb02",
  1127 => x"49c787db",
  1128 => x"c187c0fd",
  1129 => x"e2c287de",
  1130 => x"c102bfe4",
  1131 => x"c14887cb",
  1132 => x"e8e2c288",
  1133 => x"87c1c158",
  1134 => x"bfe8e2c2",
  1135 => x"87f9c002",
  1136 => x"bfe4e2c2",
  1137 => x"c280c148",
  1138 => x"c058e8e2",
  1139 => x"e2c287eb",
  1140 => x"c649bfe4",
  1141 => x"e8e2c289",
  1142 => x"a9b7c059",
  1143 => x"c287da03",
  1144 => x"c048e4e2",
  1145 => x"c287d278",
  1146 => x"02bfe8e2",
  1147 => x"e2c287cb",
  1148 => x"c648bfe4",
  1149 => x"e8e2c280",
  1150 => x"d149c058",
  1151 => x"497387dd",
  1152 => x"87e2f4c0",
  1153 => x"0e87cef1",
  1154 => x"0e5c5b5e",
  1155 => x"66cc4c71",
  1156 => x"cb4b741e",
  1157 => x"efdcc193",
  1158 => x"4aa3c483",
  1159 => x"fafe496a",
  1160 => x"c2c187d6",
  1161 => x"a3c87be2",
  1162 => x"5166d449",
  1163 => x"d849a3c9",
  1164 => x"a3ca5166",
  1165 => x"5166dc49",
  1166 => x"87d7f026",
  1167 => x"5c5b5e0e",
  1168 => x"d0ff0e5d",
  1169 => x"59a6d886",
  1170 => x"c048a6c4",
  1171 => x"c180c478",
  1172 => x"c47866c4",
  1173 => x"c478c180",
  1174 => x"c278c180",
  1175 => x"c148e8e2",
  1176 => x"cce2c278",
  1177 => x"a8de48bf",
  1178 => x"f387cb05",
  1179 => x"497087e6",
  1180 => x"ce59a6c8",
  1181 => x"e9e487ed",
  1182 => x"87cbe587",
  1183 => x"7087d8e4",
  1184 => x"acfbc04c",
  1185 => x"87d0c102",
  1186 => x"c10566d4",
  1187 => x"1ec087c2",
  1188 => x"c11ec11e",
  1189 => x"c01ed2de",
  1190 => x"87ebfd49",
  1191 => x"4a66d0c1",
  1192 => x"496a82c4",
  1193 => x"517481c7",
  1194 => x"1ed81ec1",
  1195 => x"81c8496a",
  1196 => x"d887e8e4",
  1197 => x"66c4c186",
  1198 => x"01a8c048",
  1199 => x"a6c487c7",
  1200 => x"ce78c148",
  1201 => x"66c4c187",
  1202 => x"cc88c148",
  1203 => x"87c358a6",
  1204 => x"cc87f4e3",
  1205 => x"78c248a6",
  1206 => x"cd029c74",
  1207 => x"66c487c1",
  1208 => x"66c8c148",
  1209 => x"f6cc03a8",
  1210 => x"48a6d887",
  1211 => x"80c478c0",
  1212 => x"e2e278c0",
  1213 => x"c14c7087",
  1214 => x"c205acd0",
  1215 => x"66dc87d7",
  1216 => x"87c6e57e",
  1217 => x"e0c04970",
  1218 => x"cae259a6",
  1219 => x"c04c7087",
  1220 => x"c105acec",
  1221 => x"66c487ea",
  1222 => x"c191cb49",
  1223 => x"c48166c0",
  1224 => x"4d6a4aa1",
  1225 => x"dc4aa1c8",
  1226 => x"c3c15266",
  1227 => x"e6e179e3",
  1228 => x"9c4c7087",
  1229 => x"c087d802",
  1230 => x"d202acfb",
  1231 => x"e1557487",
  1232 => x"4c7087d5",
  1233 => x"87c7029c",
  1234 => x"05acfbc0",
  1235 => x"c087eeff",
  1236 => x"c1c255e0",
  1237 => x"7d97c055",
  1238 => x"6e4966d4",
  1239 => x"87db05a9",
  1240 => x"c84866c4",
  1241 => x"ca04a866",
  1242 => x"4866c487",
  1243 => x"a6c880c1",
  1244 => x"c887c858",
  1245 => x"88c14866",
  1246 => x"e058a6cc",
  1247 => x"4c7087d9",
  1248 => x"05acd0c1",
  1249 => x"66d087c8",
  1250 => x"d480c148",
  1251 => x"d0c158a6",
  1252 => x"e9fd02ac",
  1253 => x"a6e0c087",
  1254 => x"7866d448",
  1255 => x"c04866dc",
  1256 => x"05a866e0",
  1257 => x"c087cac9",
  1258 => x"c048a6e4",
  1259 => x"48747e78",
  1260 => x"c088fbc0",
  1261 => x"7058a6ec",
  1262 => x"cfc80298",
  1263 => x"88cb4887",
  1264 => x"58a6ecc0",
  1265 => x"c1029870",
  1266 => x"c94887d2",
  1267 => x"a6ecc088",
  1268 => x"02987058",
  1269 => x"4887dbc3",
  1270 => x"ecc088c4",
  1271 => x"987058a6",
  1272 => x"4887d002",
  1273 => x"ecc088c1",
  1274 => x"987058a6",
  1275 => x"87c2c302",
  1276 => x"d887d3c7",
  1277 => x"f0c048a6",
  1278 => x"dadeff78",
  1279 => x"c04c7087",
  1280 => x"c002acec",
  1281 => x"a6dc87c3",
  1282 => x"acecc05c",
  1283 => x"ff87cd02",
  1284 => x"7087c4de",
  1285 => x"acecc04c",
  1286 => x"87f3ff05",
  1287 => x"02acecc0",
  1288 => x"ff87c4c0",
  1289 => x"d887f0dd",
  1290 => x"66d41e66",
  1291 => x"66d41e49",
  1292 => x"dec11e49",
  1293 => x"66d41ed2",
  1294 => x"87cbf749",
  1295 => x"1eca1ec0",
  1296 => x"cb4966dc",
  1297 => x"66d8c191",
  1298 => x"48a6d881",
  1299 => x"d878a1c4",
  1300 => x"ff49bf66",
  1301 => x"d887c4de",
  1302 => x"a8b7c086",
  1303 => x"87c5c106",
  1304 => x"1ede1ec1",
  1305 => x"49bf66c8",
  1306 => x"87efddff",
  1307 => x"497086c8",
  1308 => x"8808c048",
  1309 => x"c058a6dc",
  1310 => x"c006a8b7",
  1311 => x"66d887e7",
  1312 => x"a8b7dd48",
  1313 => x"6e87de03",
  1314 => x"66d849bf",
  1315 => x"51e0c081",
  1316 => x"c14966d8",
  1317 => x"81bf6e81",
  1318 => x"d851c1c2",
  1319 => x"81c24966",
  1320 => x"c081bf6e",
  1321 => x"4866cc51",
  1322 => x"a6d080c1",
  1323 => x"c47ec158",
  1324 => x"deff87da",
  1325 => x"a6dc87d4",
  1326 => x"cddeff58",
  1327 => x"a6ecc087",
  1328 => x"a8ecc058",
  1329 => x"87cac005",
  1330 => x"48a6e8c0",
  1331 => x"c07866d8",
  1332 => x"dbff87c4",
  1333 => x"66c487c1",
  1334 => x"c191cb49",
  1335 => x"714866c0",
  1336 => x"6e7e7080",
  1337 => x"6e82c84a",
  1338 => x"d881ca49",
  1339 => x"e8c05166",
  1340 => x"81c14966",
  1341 => x"c18966d8",
  1342 => x"70307148",
  1343 => x"7189c149",
  1344 => x"e6c27a97",
  1345 => x"d849bfd4",
  1346 => x"6a972966",
  1347 => x"9871484a",
  1348 => x"58a6f0c0",
  1349 => x"81c4496e",
  1350 => x"e0c04d69",
  1351 => x"66dc4866",
  1352 => x"c8c002a8",
  1353 => x"48a6d887",
  1354 => x"c5c078c0",
  1355 => x"48a6d887",
  1356 => x"66d878c1",
  1357 => x"1ee0c01e",
  1358 => x"daff4975",
  1359 => x"86c887dd",
  1360 => x"b7c04c70",
  1361 => x"d4c106ac",
  1362 => x"c0857487",
  1363 => x"897449e0",
  1364 => x"d9c14b75",
  1365 => x"fe714ad8",
  1366 => x"c287cded",
  1367 => x"66e4c085",
  1368 => x"c080c148",
  1369 => x"c058a6e8",
  1370 => x"c14966ec",
  1371 => x"02a97081",
  1372 => x"d887c8c0",
  1373 => x"78c048a6",
  1374 => x"d887c5c0",
  1375 => x"78c148a6",
  1376 => x"c21e66d8",
  1377 => x"e0c049a4",
  1378 => x"70887148",
  1379 => x"49751e49",
  1380 => x"87c7d9ff",
  1381 => x"b7c086c8",
  1382 => x"c0ff01a8",
  1383 => x"66e4c087",
  1384 => x"87d1c002",
  1385 => x"81c9496e",
  1386 => x"5166e4c0",
  1387 => x"c4c1486e",
  1388 => x"ccc078f3",
  1389 => x"c9496e87",
  1390 => x"6e51c281",
  1391 => x"e7c5c148",
  1392 => x"c07ec178",
  1393 => x"d7ff87c6",
  1394 => x"4c7087fd",
  1395 => x"f5c0026e",
  1396 => x"4866c487",
  1397 => x"04a866c8",
  1398 => x"c487cbc0",
  1399 => x"80c14866",
  1400 => x"c058a6c8",
  1401 => x"66c887e0",
  1402 => x"cc88c148",
  1403 => x"d5c058a6",
  1404 => x"acc6c187",
  1405 => x"87c8c005",
  1406 => x"c14866cc",
  1407 => x"58a6d080",
  1408 => x"87c3d7ff",
  1409 => x"66d04c70",
  1410 => x"d480c148",
  1411 => x"9c7458a6",
  1412 => x"87cbc002",
  1413 => x"c14866c4",
  1414 => x"04a866c8",
  1415 => x"ff87caf3",
  1416 => x"c487dbd6",
  1417 => x"a8c74866",
  1418 => x"87e5c003",
  1419 => x"48e8e2c2",
  1420 => x"66c478c0",
  1421 => x"c191cb49",
  1422 => x"c48166c0",
  1423 => x"4a6a4aa1",
  1424 => x"c47952c0",
  1425 => x"80c14866",
  1426 => x"c758a6c8",
  1427 => x"dbff04a8",
  1428 => x"8ed0ff87",
  1429 => x"87f9dfff",
  1430 => x"1e00203a",
  1431 => x"4b711e73",
  1432 => x"87c6029b",
  1433 => x"48e4e2c2",
  1434 => x"1ec778c0",
  1435 => x"bfe4e2c2",
  1436 => x"dcc11e49",
  1437 => x"e2c21eef",
  1438 => x"ee49bfcc",
  1439 => x"86cc87fe",
  1440 => x"bfcce2c2",
  1441 => x"87c3ea49",
  1442 => x"c8029b73",
  1443 => x"efdcc187",
  1444 => x"e3e3c049",
  1445 => x"fcdeff87",
  1446 => x"d4c71e87",
  1447 => x"fe49c187",
  1448 => x"f0fe87f9",
  1449 => x"987087d0",
  1450 => x"fe87cd02",
  1451 => x"7087e9f7",
  1452 => x"87c40298",
  1453 => x"87c24ac1",
  1454 => x"9a724ac0",
  1455 => x"c087ce05",
  1456 => x"eadbc11e",
  1457 => x"faf0c049",
  1458 => x"fe86c487",
  1459 => x"c11ec087",
  1460 => x"c049f5db",
  1461 => x"c087ecf0",
  1462 => x"d5f6c01e",
  1463 => x"c0497087",
  1464 => x"c387e0f0",
  1465 => x"8ef887ca",
  1466 => x"44534f26",
  1467 => x"69616620",
  1468 => x"2e64656c",
  1469 => x"6f6f4200",
  1470 => x"676e6974",
  1471 => x"002e2e2e",
  1472 => x"d4e7c01e",
  1473 => x"2687fa87",
  1474 => x"e2c21e4f",
  1475 => x"78c048e4",
  1476 => x"48cce2c2",
  1477 => x"c0fe78c0",
  1478 => x"c087e587",
  1479 => x"004f2648",
  1480 => x"45208000",
  1481 => x"00746978",
  1482 => x"61422080",
  1483 => x"e3006b63",
  1484 => x"b8000010",
  1485 => x"00000028",
  1486 => x"10e30000",
  1487 => x"28d60000",
  1488 => x"00000000",
  1489 => x"0010e300",
  1490 => x"0028f400",
  1491 => x"00000000",
  1492 => x"000010e3",
  1493 => x"00002912",
  1494 => x"e3000000",
  1495 => x"30000010",
  1496 => x"00000029",
  1497 => x"10e30000",
  1498 => x"294e0000",
  1499 => x"00000000",
  1500 => x"0010e300",
  1501 => x"00296c00",
  1502 => x"00000000",
  1503 => x"000010e3",
  1504 => x"00000000",
  1505 => x"78000000",
  1506 => x"00000011",
  1507 => x"00000000",
  1508 => x"6f4c0000",
  1509 => x"2a206461",
  1510 => x"fe1e002e",
  1511 => x"78c048f0",
  1512 => x"097909cd",
  1513 => x"1e1e4f26",
  1514 => x"7ebff0fe",
  1515 => x"4f262648",
  1516 => x"48f0fe1e",
  1517 => x"4f2678c1",
  1518 => x"48f0fe1e",
  1519 => x"4f2678c0",
  1520 => x"c04a711e",
  1521 => x"4f265252",
  1522 => x"5c5b5e0e",
  1523 => x"86f40e5d",
  1524 => x"6d974d71",
  1525 => x"4ca5c17e",
  1526 => x"c8486c97",
  1527 => x"486e58a6",
  1528 => x"05a866c4",
  1529 => x"48ff87c5",
  1530 => x"ff87e6c0",
  1531 => x"a5c287ca",
  1532 => x"4b6c9749",
  1533 => x"974ba371",
  1534 => x"6c974b6b",
  1535 => x"c1486e7e",
  1536 => x"58a6c880",
  1537 => x"a6cc98c7",
  1538 => x"7c977058",
  1539 => x"7387e1fe",
  1540 => x"268ef448",
  1541 => x"264c264d",
  1542 => x"0e4f264b",
  1543 => x"0e5c5b5e",
  1544 => x"4c7186f4",
  1545 => x"c34a66d8",
  1546 => x"a4c29aff",
  1547 => x"496c974b",
  1548 => x"7249a173",
  1549 => x"7e6c9751",
  1550 => x"80c1486e",
  1551 => x"c758a6c8",
  1552 => x"58a6cc98",
  1553 => x"8ef45470",
  1554 => x"1e87caff",
  1555 => x"87e8fd1e",
  1556 => x"494abfe0",
  1557 => x"99c0e0c0",
  1558 => x"7287cb02",
  1559 => x"cae6c21e",
  1560 => x"87f7fe49",
  1561 => x"fdfc86c4",
  1562 => x"fd7e7087",
  1563 => x"262687c2",
  1564 => x"e6c21e4f",
  1565 => x"c7fd49ca",
  1566 => x"cbe1c187",
  1567 => x"87dafc49",
  1568 => x"2687dcc3",
  1569 => x"4f261e4f",
  1570 => x"5c5b5e0e",
  1571 => x"c24c710e",
  1572 => x"fc49cae6",
  1573 => x"4a7087f2",
  1574 => x"04aab7c0",
  1575 => x"c387e3c2",
  1576 => x"c905aae0",
  1577 => x"d2e5c187",
  1578 => x"c278c148",
  1579 => x"f0c387d4",
  1580 => x"87c905aa",
  1581 => x"48cee5c1",
  1582 => x"f5c178c1",
  1583 => x"d2e5c187",
  1584 => x"87c702bf",
  1585 => x"c0c24b72",
  1586 => x"7287c2b3",
  1587 => x"059c744b",
  1588 => x"e5c187d1",
  1589 => x"c11ebfce",
  1590 => x"1ebfd2e5",
  1591 => x"e4fe4972",
  1592 => x"c186c887",
  1593 => x"02bfcee5",
  1594 => x"7387e0c0",
  1595 => x"29b7c449",
  1596 => x"eee6c191",
  1597 => x"cf4a7381",
  1598 => x"c192c29a",
  1599 => x"70307248",
  1600 => x"72baff4a",
  1601 => x"70986948",
  1602 => x"7387db79",
  1603 => x"29b7c449",
  1604 => x"eee6c191",
  1605 => x"cf4a7381",
  1606 => x"c392c29a",
  1607 => x"70307248",
  1608 => x"b069484a",
  1609 => x"e5c17970",
  1610 => x"78c048d2",
  1611 => x"48cee5c1",
  1612 => x"e6c278c0",
  1613 => x"cffa49ca",
  1614 => x"c04a7087",
  1615 => x"fd03aab7",
  1616 => x"48c087dd",
  1617 => x"4d2687c2",
  1618 => x"4b264c26",
  1619 => x"00004f26",
  1620 => x"00000000",
  1621 => x"711e0000",
  1622 => x"ebfc494a",
  1623 => x"1e4f2687",
  1624 => x"49724ac0",
  1625 => x"e6c191c4",
  1626 => x"79c081ee",
  1627 => x"b7d082c1",
  1628 => x"87ee04aa",
  1629 => x"5e0e4f26",
  1630 => x"0e5d5c5b",
  1631 => x"f7f84d71",
  1632 => x"c44a7587",
  1633 => x"c1922ab7",
  1634 => x"7582eee6",
  1635 => x"c29ccf4c",
  1636 => x"4b496a94",
  1637 => x"9bc32b74",
  1638 => x"307448c2",
  1639 => x"bcff4c70",
  1640 => x"98714874",
  1641 => x"c7f87a70",
  1642 => x"fe487387",
  1643 => x"000087d8",
  1644 => x"00000000",
  1645 => x"00000000",
  1646 => x"00000000",
  1647 => x"00000000",
  1648 => x"00000000",
  1649 => x"00000000",
  1650 => x"00000000",
  1651 => x"00000000",
  1652 => x"00000000",
  1653 => x"00000000",
  1654 => x"00000000",
  1655 => x"00000000",
  1656 => x"00000000",
  1657 => x"00000000",
  1658 => x"00000000",
  1659 => x"ff1e0000",
  1660 => x"e1c848d0",
  1661 => x"ff487178",
  1662 => x"c47808d4",
  1663 => x"d4ff4866",
  1664 => x"4f267808",
  1665 => x"c44a711e",
  1666 => x"721e4966",
  1667 => x"87deff49",
  1668 => x"c048d0ff",
  1669 => x"262678e0",
  1670 => x"1e731e4f",
  1671 => x"66c84b71",
  1672 => x"4a731e49",
  1673 => x"49a2e0c1",
  1674 => x"2687d9ff",
  1675 => x"4d2687c4",
  1676 => x"4b264c26",
  1677 => x"711e4f26",
  1678 => x"da1e494a",
  1679 => x"87eefe49",
  1680 => x"49bf66c8",
  1681 => x"c44866c8",
  1682 => x"58a6cc80",
  1683 => x"ff29b7c8",
  1684 => x"787148d4",
  1685 => x"49bf66c8",
  1686 => x"7129b7c8",
  1687 => x"48d0ff78",
  1688 => x"2678e0c0",
  1689 => x"ff1e4f26",
  1690 => x"ffc34ad4",
  1691 => x"48d0ff7a",
  1692 => x"de78e1c0",
  1693 => x"d4e6c27a",
  1694 => x"48497abf",
  1695 => x"7a7028c8",
  1696 => x"28d04871",
  1697 => x"48717a70",
  1698 => x"7a7028d8",
  1699 => x"c048d0ff",
  1700 => x"4f2678e0",
  1701 => x"5c5b5e0e",
  1702 => x"4c710e5d",
  1703 => x"bfd4e6c2",
  1704 => x"2b744b4d",
  1705 => x"c19b66d0",
  1706 => x"ab66d483",
  1707 => x"c087c204",
  1708 => x"d04a744b",
  1709 => x"31724966",
  1710 => x"9975b9ff",
  1711 => x"30724873",
  1712 => x"71484a70",
  1713 => x"d8e6c2b0",
  1714 => x"87dafe58",
  1715 => x"4c264d26",
  1716 => x"4f264b26",
  1717 => x"48d0ff1e",
  1718 => x"7178c9c8",
  1719 => x"08d4ff48",
  1720 => x"1e4f2678",
  1721 => x"eb494a71",
  1722 => x"48d0ff87",
  1723 => x"4f2678c8",
  1724 => x"711e731e",
  1725 => x"e4e6c24b",
  1726 => x"87c302bf",
  1727 => x"ff87ebc2",
  1728 => x"c9c848d0",
  1729 => x"c0497378",
  1730 => x"d4ffb1e0",
  1731 => x"c2787148",
  1732 => x"c048d8e6",
  1733 => x"0266c878",
  1734 => x"ffc387c5",
  1735 => x"c087c249",
  1736 => x"e0e6c249",
  1737 => x"0266cc59",
  1738 => x"d5c587c6",
  1739 => x"87c44ad5",
  1740 => x"4affffcf",
  1741 => x"5ae4e6c2",
  1742 => x"48e4e6c2",
  1743 => x"87c478c1",
  1744 => x"4c264d26",
  1745 => x"4f264b26",
  1746 => x"5c5b5e0e",
  1747 => x"4a710e5d",
  1748 => x"bfe0e6c2",
  1749 => x"029a724c",
  1750 => x"c84987cb",
  1751 => x"e6ebc191",
  1752 => x"c483714b",
  1753 => x"e6efc187",
  1754 => x"134dc04b",
  1755 => x"c2997449",
  1756 => x"b9bfdce6",
  1757 => x"7148d4ff",
  1758 => x"2cb7c178",
  1759 => x"adb7c885",
  1760 => x"c287e804",
  1761 => x"48bfd8e6",
  1762 => x"e6c280c8",
  1763 => x"effe58dc",
  1764 => x"1e731e87",
  1765 => x"4a134b71",
  1766 => x"87cb029a",
  1767 => x"e7fe4972",
  1768 => x"9a4a1387",
  1769 => x"fe87f505",
  1770 => x"c21e87da",
  1771 => x"49bfd8e6",
  1772 => x"48d8e6c2",
  1773 => x"c478a1c1",
  1774 => x"03a9b7c0",
  1775 => x"d4ff87db",
  1776 => x"dce6c248",
  1777 => x"e6c278bf",
  1778 => x"c249bfd8",
  1779 => x"c148d8e6",
  1780 => x"c0c478a1",
  1781 => x"e504a9b7",
  1782 => x"48d0ff87",
  1783 => x"e6c278c8",
  1784 => x"78c048e4",
  1785 => x"00004f26",
  1786 => x"00000000",
  1787 => x"00000000",
  1788 => x"005f5f00",
  1789 => x"03000000",
  1790 => x"03030003",
  1791 => x"7f140000",
  1792 => x"7f7f147f",
  1793 => x"24000014",
  1794 => x"3a6b6b2e",
  1795 => x"6a4c0012",
  1796 => x"566c1836",
  1797 => x"7e300032",
  1798 => x"3a77594f",
  1799 => x"00004068",
  1800 => x"00030704",
  1801 => x"00000000",
  1802 => x"41633e1c",
  1803 => x"00000000",
  1804 => x"1c3e6341",
  1805 => x"2a080000",
  1806 => x"3e1c1c3e",
  1807 => x"0800082a",
  1808 => x"083e3e08",
  1809 => x"00000008",
  1810 => x"0060e080",
  1811 => x"08000000",
  1812 => x"08080808",
  1813 => x"00000008",
  1814 => x"00606000",
  1815 => x"60400000",
  1816 => x"060c1830",
  1817 => x"3e000103",
  1818 => x"7f4d597f",
  1819 => x"0400003e",
  1820 => x"007f7f06",
  1821 => x"42000000",
  1822 => x"4f597163",
  1823 => x"22000046",
  1824 => x"7f494963",
  1825 => x"1c180036",
  1826 => x"7f7f1316",
  1827 => x"27000010",
  1828 => x"7d454567",
  1829 => x"3c000039",
  1830 => x"79494b7e",
  1831 => x"01000030",
  1832 => x"0f797101",
  1833 => x"36000007",
  1834 => x"7f49497f",
  1835 => x"06000036",
  1836 => x"3f69494f",
  1837 => x"0000001e",
  1838 => x"00666600",
  1839 => x"00000000",
  1840 => x"0066e680",
  1841 => x"08000000",
  1842 => x"22141408",
  1843 => x"14000022",
  1844 => x"14141414",
  1845 => x"22000014",
  1846 => x"08141422",
  1847 => x"02000008",
  1848 => x"0f595103",
  1849 => x"7f3e0006",
  1850 => x"1f555d41",
  1851 => x"7e00001e",
  1852 => x"7f09097f",
  1853 => x"7f00007e",
  1854 => x"7f49497f",
  1855 => x"1c000036",
  1856 => x"4141633e",
  1857 => x"7f000041",
  1858 => x"3e63417f",
  1859 => x"7f00001c",
  1860 => x"4149497f",
  1861 => x"7f000041",
  1862 => x"0109097f",
  1863 => x"3e000001",
  1864 => x"7b49417f",
  1865 => x"7f00007a",
  1866 => x"7f08087f",
  1867 => x"0000007f",
  1868 => x"417f7f41",
  1869 => x"20000000",
  1870 => x"7f404060",
  1871 => x"7f7f003f",
  1872 => x"63361c08",
  1873 => x"7f000041",
  1874 => x"4040407f",
  1875 => x"7f7f0040",
  1876 => x"7f060c06",
  1877 => x"7f7f007f",
  1878 => x"7f180c06",
  1879 => x"3e00007f",
  1880 => x"7f41417f",
  1881 => x"7f00003e",
  1882 => x"0f09097f",
  1883 => x"7f3e0006",
  1884 => x"7e7f6141",
  1885 => x"7f000040",
  1886 => x"7f19097f",
  1887 => x"26000066",
  1888 => x"7b594d6f",
  1889 => x"01000032",
  1890 => x"017f7f01",
  1891 => x"3f000001",
  1892 => x"7f40407f",
  1893 => x"0f00003f",
  1894 => x"3f70703f",
  1895 => x"7f7f000f",
  1896 => x"7f301830",
  1897 => x"6341007f",
  1898 => x"361c1c36",
  1899 => x"03014163",
  1900 => x"067c7c06",
  1901 => x"71610103",
  1902 => x"43474d59",
  1903 => x"00000041",
  1904 => x"41417f7f",
  1905 => x"03010000",
  1906 => x"30180c06",
  1907 => x"00004060",
  1908 => x"7f7f4141",
  1909 => x"0c080000",
  1910 => x"0c060306",
  1911 => x"80800008",
  1912 => x"80808080",
  1913 => x"00000080",
  1914 => x"04070300",
  1915 => x"20000000",
  1916 => x"7c545474",
  1917 => x"7f000078",
  1918 => x"7c44447f",
  1919 => x"38000038",
  1920 => x"4444447c",
  1921 => x"38000000",
  1922 => x"7f44447c",
  1923 => x"3800007f",
  1924 => x"5c54547c",
  1925 => x"04000018",
  1926 => x"05057f7e",
  1927 => x"18000000",
  1928 => x"fca4a4bc",
  1929 => x"7f00007c",
  1930 => x"7c04047f",
  1931 => x"00000078",
  1932 => x"407d3d00",
  1933 => x"80000000",
  1934 => x"7dfd8080",
  1935 => x"7f000000",
  1936 => x"6c38107f",
  1937 => x"00000044",
  1938 => x"407f3f00",
  1939 => x"7c7c0000",
  1940 => x"7c0c180c",
  1941 => x"7c000078",
  1942 => x"7c04047c",
  1943 => x"38000078",
  1944 => x"7c44447c",
  1945 => x"fc000038",
  1946 => x"3c2424fc",
  1947 => x"18000018",
  1948 => x"fc24243c",
  1949 => x"7c0000fc",
  1950 => x"0c04047c",
  1951 => x"48000008",
  1952 => x"7454545c",
  1953 => x"04000020",
  1954 => x"44447f3f",
  1955 => x"3c000000",
  1956 => x"7c40407c",
  1957 => x"1c00007c",
  1958 => x"3c60603c",
  1959 => x"7c3c001c",
  1960 => x"7c603060",
  1961 => x"6c44003c",
  1962 => x"6c381038",
  1963 => x"1c000044",
  1964 => x"3c60e0bc",
  1965 => x"4400001c",
  1966 => x"4c5c7464",
  1967 => x"08000044",
  1968 => x"41773e08",
  1969 => x"00000041",
  1970 => x"007f7f00",
  1971 => x"41000000",
  1972 => x"083e7741",
  1973 => x"01020008",
  1974 => x"02020301",
  1975 => x"7f7f0001",
  1976 => x"7f7f7f7f",
  1977 => x"0808007f",
  1978 => x"3e3e1c1c",
  1979 => x"7f7f7f7f",
  1980 => x"1c1c3e3e",
  1981 => x"10000808",
  1982 => x"187c7c18",
  1983 => x"10000010",
  1984 => x"307c7c30",
  1985 => x"30100010",
  1986 => x"1e786060",
  1987 => x"66420006",
  1988 => x"663c183c",
  1989 => x"38780042",
  1990 => x"6cc6c26a",
  1991 => x"00600038",
  1992 => x"00006000",
  1993 => x"5e0e0060",
  1994 => x"0e5d5c5b",
  1995 => x"c24c711e",
  1996 => x"4dbff5e6",
  1997 => x"1ec04bc0",
  1998 => x"c702ab74",
  1999 => x"48a6c487",
  2000 => x"87c578c0",
  2001 => x"c148a6c4",
  2002 => x"1e66c478",
  2003 => x"dfee4973",
  2004 => x"c086c887",
  2005 => x"efef49e0",
  2006 => x"4aa5c487",
  2007 => x"f0f0496a",
  2008 => x"87c6f187",
  2009 => x"83c185cb",
  2010 => x"04abb7c8",
  2011 => x"2687c7ff",
  2012 => x"4c264d26",
  2013 => x"4f264b26",
  2014 => x"c24a711e",
  2015 => x"c25af9e6",
  2016 => x"c748f9e6",
  2017 => x"ddfe4978",
  2018 => x"1e4f2687",
  2019 => x"4a711e73",
  2020 => x"03aab7c0",
  2021 => x"cdc287d3",
  2022 => x"c405bfd8",
  2023 => x"c24bc187",
  2024 => x"c24bc087",
  2025 => x"c45bdccd",
  2026 => x"dccdc287",
  2027 => x"d8cdc25a",
  2028 => x"9ac14abf",
  2029 => x"49a2c0c1",
  2030 => x"fc87e8ec",
  2031 => x"d8cdc248",
  2032 => x"effe78bf",
  2033 => x"5b5e0e87",
  2034 => x"710e5d5c",
  2035 => x"f84a6b4b",
  2036 => x"c74dc0c4",
  2037 => x"d04cc0fc",
  2038 => x"99c24966",
  2039 => x"d487cf02",
  2040 => x"09c04966",
  2041 => x"c84c7189",
  2042 => x"8a66d434",
  2043 => x"66d087d7",
  2044 => x"0299c149",
  2045 => x"66d487ca",
  2046 => x"d435c84d",
  2047 => x"87c58266",
  2048 => x"b7c492cf",
  2049 => x"aab7752a",
  2050 => x"4a87c103",
  2051 => x"06aab774",
  2052 => x"724a87c1",
  2053 => x"87d8fd7b",
  2054 => x"d8cdc21e",
  2055 => x"f5e449bf",
  2056 => x"ede6c287",
  2057 => x"78bfe848",
  2058 => x"48e9e6c2",
  2059 => x"c278bfec",
  2060 => x"4abfede6",
  2061 => x"99ffc349",
  2062 => x"722ab7c8",
  2063 => x"c2b07148",
  2064 => x"2658f5e6",
  2065 => x"5b5e0e4f",
  2066 => x"710e5d5c",
  2067 => x"87c8ff4b",
  2068 => x"48e8e6c2",
  2069 => x"497350c0",
  2070 => x"7087dbe4",
  2071 => x"9cc24c49",
  2072 => x"cb49eecb",
  2073 => x"497087fa",
  2074 => x"e8e6c24d",
  2075 => x"c105bf97",
  2076 => x"66d087e2",
  2077 => x"f1e6c249",
  2078 => x"d60599bf",
  2079 => x"4966d487",
  2080 => x"bfe9e6c2",
  2081 => x"87cb0599",
  2082 => x"e9e34973",
  2083 => x"02987087",
  2084 => x"c187c1c1",
  2085 => x"87c0fe4c",
  2086 => x"cfcb4975",
  2087 => x"02987087",
  2088 => x"e6c287c6",
  2089 => x"50c148e8",
  2090 => x"97e8e6c2",
  2091 => x"e3c005bf",
  2092 => x"f1e6c287",
  2093 => x"66d049bf",
  2094 => x"d6ff0599",
  2095 => x"e9e6c287",
  2096 => x"66d449bf",
  2097 => x"caff0599",
  2098 => x"e2497387",
  2099 => x"987087e8",
  2100 => x"87fffe05",
  2101 => x"d7fa4874",
  2102 => x"5b5e0e87",
  2103 => x"f40e5d5c",
  2104 => x"4c4dc086",
  2105 => x"c47ebfec",
  2106 => x"e6c248a6",
  2107 => x"c178bff5",
  2108 => x"c71ec01e",
  2109 => x"87cdfd49",
  2110 => x"987086c8",
  2111 => x"ff87cd02",
  2112 => x"87c7fa49",
  2113 => x"e149dac1",
  2114 => x"4dc187ec",
  2115 => x"97e8e6c2",
  2116 => x"87c302bf",
  2117 => x"c287eec9",
  2118 => x"4bbfede6",
  2119 => x"bfd8cdc2",
  2120 => x"87d9c105",
  2121 => x"c848a6c4",
  2122 => x"c278c0c0",
  2123 => x"6e7eddd4",
  2124 => x"6e49bf97",
  2125 => x"7080c148",
  2126 => x"f9e0717e",
  2127 => x"02987087",
  2128 => x"66c487c3",
  2129 => x"4866c4b3",
  2130 => x"c828b7c1",
  2131 => x"987058a6",
  2132 => x"87dbff05",
  2133 => x"e049fdc3",
  2134 => x"fac387dc",
  2135 => x"87d6e049",
  2136 => x"ffc34973",
  2137 => x"c01e7199",
  2138 => x"87c6c949",
  2139 => x"b7c84973",
  2140 => x"c11e7129",
  2141 => x"87fac849",
  2142 => x"c1c686c8",
  2143 => x"f1e6c287",
  2144 => x"029b4bbf",
  2145 => x"cdc287dd",
  2146 => x"c749bfd4",
  2147 => x"987087de",
  2148 => x"c087c405",
  2149 => x"c287d24b",
  2150 => x"c3c749e0",
  2151 => x"d8cdc287",
  2152 => x"c287c658",
  2153 => x"c048d4cd",
  2154 => x"c2497378",
  2155 => x"87ce0599",
  2156 => x"ff49ebc3",
  2157 => x"7087ffde",
  2158 => x"0299c249",
  2159 => x"4cfb87c2",
  2160 => x"99c14973",
  2161 => x"c387ce05",
  2162 => x"deff49f4",
  2163 => x"497087e8",
  2164 => x"c20299c2",
  2165 => x"734cfa87",
  2166 => x"0599c849",
  2167 => x"f5c387ce",
  2168 => x"d1deff49",
  2169 => x"c2497087",
  2170 => x"87d50299",
  2171 => x"bff9e6c2",
  2172 => x"4887ca02",
  2173 => x"e6c288c1",
  2174 => x"c2c058fd",
  2175 => x"c14cff87",
  2176 => x"c449734d",
  2177 => x"87ce0599",
  2178 => x"ff49f2c3",
  2179 => x"7087e7dd",
  2180 => x"0299c249",
  2181 => x"e6c287dc",
  2182 => x"487ebff9",
  2183 => x"03a8b7c7",
  2184 => x"6e87cbc0",
  2185 => x"c280c148",
  2186 => x"c058fde6",
  2187 => x"4cfe87c2",
  2188 => x"fdc34dc1",
  2189 => x"fddcff49",
  2190 => x"c2497087",
  2191 => x"d5c00299",
  2192 => x"f9e6c287",
  2193 => x"c9c002bf",
  2194 => x"f9e6c287",
  2195 => x"c078c048",
  2196 => x"4cfd87c2",
  2197 => x"fac34dc1",
  2198 => x"d9dcff49",
  2199 => x"c2497087",
  2200 => x"d9c00299",
  2201 => x"f9e6c287",
  2202 => x"b7c748bf",
  2203 => x"c9c003a8",
  2204 => x"f9e6c287",
  2205 => x"c078c748",
  2206 => x"4cfc87c2",
  2207 => x"b7c04dc1",
  2208 => x"d1c003ac",
  2209 => x"4a66c487",
  2210 => x"6a82d8c1",
  2211 => x"87c6c002",
  2212 => x"49744b6a",
  2213 => x"1ec00f73",
  2214 => x"c11ef0c3",
  2215 => x"e4f649da",
  2216 => x"7086c887",
  2217 => x"e2c00298",
  2218 => x"48a6c887",
  2219 => x"bff9e6c2",
  2220 => x"4966c878",
  2221 => x"66c491cb",
  2222 => x"70807148",
  2223 => x"02bf6e7e",
  2224 => x"6e87c8c0",
  2225 => x"66c84bbf",
  2226 => x"750f7349",
  2227 => x"c8c0029d",
  2228 => x"f9e6c287",
  2229 => x"cdf149bf",
  2230 => x"dccdc287",
  2231 => x"ddc002bf",
  2232 => x"c7c24987",
  2233 => x"02987087",
  2234 => x"c287d3c0",
  2235 => x"49bff9e6",
  2236 => x"c087f3f0",
  2237 => x"87d3f249",
  2238 => x"48dccdc2",
  2239 => x"8ef478c0",
  2240 => x"0e87edf1",
  2241 => x"5d5c5b5e",
  2242 => x"4c711e0e",
  2243 => x"bff5e6c2",
  2244 => x"a1cdc149",
  2245 => x"81d1c14d",
  2246 => x"9c747e69",
  2247 => x"c487cf02",
  2248 => x"7b744ba5",
  2249 => x"bff5e6c2",
  2250 => x"87ccf149",
  2251 => x"9c747b6e",
  2252 => x"c087c405",
  2253 => x"c187c24b",
  2254 => x"f149734b",
  2255 => x"66d487cd",
  2256 => x"4987c702",
  2257 => x"4a7087da",
  2258 => x"4ac087c2",
  2259 => x"5ae0cdc2",
  2260 => x"87dcf026",
  2261 => x"00000000",
  2262 => x"00000000",
  2263 => x"00000000",
  2264 => x"ff4a711e",
  2265 => x"7249bfc8",
  2266 => x"4f2648a1",
  2267 => x"bfc8ff1e",
  2268 => x"c0c0fe89",
  2269 => x"a9c0c0c0",
  2270 => x"c087c401",
  2271 => x"c187c24a",
  2272 => x"2648724a",
  2273 => x"cec21e4f",
  2274 => x"c149bfee",
  2275 => x"f2cec2b9",
  2276 => x"48d4ff59",
  2277 => x"ff78ffc3",
  2278 => x"e1c048d0",
  2279 => x"48d4ff78",
  2280 => x"31c478c1",
  2281 => x"d0ff7871",
  2282 => x"78e0c048",
  2283 => x"00004f26",
  2284 => x"5e0e0000",
  2285 => x"0e5d5c5b",
  2286 => x"bfec4d71",
  2287 => x"ff49c54b",
  2288 => x"7087f3d6",
  2289 => x"87c70598",
  2290 => x"99c24973",
  2291 => x"c287c702",
  2292 => x"c248edd4",
  2293 => x"49c678c0",
  2294 => x"87dad6ff",
  2295 => x"c7059870",
  2296 => x"c4497387",
  2297 => x"87c70299",
  2298 => x"48edd4c2",
  2299 => x"c478f0c0",
  2300 => x"c1d6ff49",
  2301 => x"05987087",
  2302 => x"497387c7",
  2303 => x"c60299c8",
  2304 => x"edd4c287",
  2305 => x"cc78cc48",
  2306 => x"e9d5ff49",
  2307 => x"05987087",
  2308 => x"497387c7",
  2309 => x"c60299d0",
  2310 => x"edd4c287",
  2311 => x"d078c848",
  2312 => x"49751e66",
  2313 => x"87f1d7ff",
  2314 => x"bfedd4c2",
  2315 => x"1e66d81e",
  2316 => x"93c24b75",
  2317 => x"94c84c75",
  2318 => x"84fde6c2",
  2319 => x"c4ee496c",
  2320 => x"c27c7087",
  2321 => x"1ebfedd4",
  2322 => x"4966e0c0",
  2323 => x"7129b7c2",
  2324 => x"c293c41e",
  2325 => x"6b83c1e7",
  2326 => x"87e9ed49",
  2327 => x"e6c27b70",
  2328 => x"49751efd",
  2329 => x"87ced7ff",
  2330 => x"4d268ee8",
  2331 => x"4b264c26",
  2332 => x"731e4f26",
  2333 => x"dfdcc11e",
  2334 => x"c250c048",
  2335 => x"c248f0d4",
  2336 => x"c278c0c0",
  2337 => x"48bfd4e6",
  2338 => x"e6c2b0c1",
  2339 => x"d7ff58d8",
  2340 => x"d3c287d4",
  2341 => x"e3fe49ee",
  2342 => x"4b7087c2",
  2343 => x"bfd4e6c2",
  2344 => x"c298fe48",
  2345 => x"ff58d8e6",
  2346 => x"7387fbd6",
  2347 => x"87c7059b",
  2348 => x"48fad3c2",
  2349 => x"c287f4c0",
  2350 => x"48bfd4e6",
  2351 => x"e6c2b0c1",
  2352 => x"d6ff58d8",
  2353 => x"d4c287e0",
  2354 => x"78c148f0",
  2355 => x"48dfdcc1",
  2356 => x"d4c250c1",
  2357 => x"e2fe49d1",
  2358 => x"e6c287c2",
  2359 => x"fe48bfd4",
  2360 => x"d8e6c298",
  2361 => x"fdd5ff58",
  2362 => x"fe48c087",
  2363 => x"455687c0",
  2364 => x"45525443",
  2365 => x"49422058",
  2366 => x"4556004e",
  2367 => x"45525443",
  2368 => x"49422e58",
  2369 => x"6f6e204e",
  2370 => x"6f662074",
  2371 => x"21646e75",
  2372 => x"54554100",
  2373 => x"4f4f424f",
  2374 => x"43455654",
  2375 => x"14125800",
  2376 => x"1c1b1d11",
  2377 => x"494a5923",
  2378 => x"ebf2f541",
  2379 => x"000080f4",
  2380 => x"00008000",
  others => ( x"00000000")
);

-- Xilinx Vivado attributes
attribute ram_style: string;
attribute ram_style of ram: signal is "block";

signal q_local : std_logic_vector((NB_COL * COL_WIDTH)-1 downto 0);

signal wea : std_logic_vector(NB_COL - 1 downto 0);

begin

	output:
	for i in 0 to NB_COL - 1 generate
		q((i + 1) * COL_WIDTH - 1 downto i * COL_WIDTH) <= q_local((i+1) * COL_WIDTH - 1 downto i * COL_WIDTH);
	end generate;
    
    -- Generate write enable signals
    -- The Block ram generator doesn't like it when the compare is done in the if statement it self.
    wea <= bytesel when we = '1' else (others => '0');

    process(clk)
    begin
        if rising_edge(clk) then
            q_local <= ram(to_integer(unsigned(addr)));
            for i in 0 to NB_COL - 1 loop
                if (wea(NB_COL-i-1) = '1') then
                    ram(to_integer(unsigned(addr)))((i + 1) * COL_WIDTH - 1 downto i * COL_WIDTH) <= d((i + 1) * COL_WIDTH - 1 downto i * COL_WIDTH);
                end if;
            end loop;
        end if;
    end process;

end arch;
